module MLP_model (
    input predict,
    input [783:0] inp,
    output reg [3:0] class
);

    // Layer 1: Dense
    reg signed [5:0] layer_1_weights [783:0][15:0];
    reg signed [5:0] layer_1_biases [15:0];
    reg signed [6:0] layer_1_outputs [15:0];

    // Layer 2: Dense
    reg signed [5:0] layer_2_weights [15:0][9:0];
    reg signed [5:0] layer_2_biases [9:0];
    reg signed [13:0] layer_2_outputs [9:0];

    reg signed [13:0] max_val;
    reg [3:0] max_idx;

    initial begin
        layer_1_weights[0][0] = -1;
        layer_1_weights[1][0] = 0;
        layer_1_weights[2][0] = 0;
        layer_1_weights[3][0] = 0;
        layer_1_weights[4][0] = -1;
        layer_1_weights[5][0] = 0;
        layer_1_weights[6][0] = 0;
        layer_1_weights[7][0] = 1;
        layer_1_weights[8][0] = 0;
        layer_1_weights[9][0] = 0;
        layer_1_weights[10][0] = 0;
        layer_1_weights[11][0] = 0;
        layer_1_weights[12][0] = 1;
        layer_1_weights[13][0] = 1;
        layer_1_weights[14][0] = 0;
        layer_1_weights[15][0] = -1;
        layer_1_weights[16][0] = 0;
        layer_1_weights[17][0] = 1;
        layer_1_weights[18][0] = -1;
        layer_1_weights[19][0] = 0;
        layer_1_weights[20][0] = 0;
        layer_1_weights[21][0] = -1;
        layer_1_weights[22][0] = 0;
        layer_1_weights[23][0] = 0;
        layer_1_weights[24][0] = -1;
        layer_1_weights[25][0] = 0;
        layer_1_weights[26][0] = 0;
        layer_1_weights[27][0] = 1;
        layer_1_weights[28][0] = 0;
        layer_1_weights[29][0] = 0;
        layer_1_weights[30][0] = 0;
        layer_1_weights[31][0] = -1;
        layer_1_weights[32][0] = 0;
        layer_1_weights[33][0] = 3;
        layer_1_weights[34][0] = 3;
        layer_1_weights[35][0] = 4;
        layer_1_weights[36][0] = 3;
        layer_1_weights[37][0] = 3;
        layer_1_weights[38][0] = 3;
        layer_1_weights[39][0] = 0;
        layer_1_weights[40][0] = 3;
        layer_1_weights[41][0] = 2;
        layer_1_weights[42][0] = 0;
        layer_1_weights[43][0] = 4;
        layer_1_weights[44][0] = 3;
        layer_1_weights[45][0] = 5;
        layer_1_weights[46][0] = 5;
        layer_1_weights[47][0] = 5;
        layer_1_weights[48][0] = 4;
        layer_1_weights[49][0] = 4;
        layer_1_weights[50][0] = 3;
        layer_1_weights[51][0] = 1;
        layer_1_weights[52][0] = -1;
        layer_1_weights[53][0] = 0;
        layer_1_weights[54][0] = 0;
        layer_1_weights[55][0] = 0;
        layer_1_weights[56][0] = -1;
        layer_1_weights[57][0] = 0;
        layer_1_weights[58][0] = 1;
        layer_1_weights[59][0] = -1;
        layer_1_weights[60][0] = 3;
        layer_1_weights[61][0] = 1;
        layer_1_weights[62][0] = 3;
        layer_1_weights[63][0] = 4;
        layer_1_weights[64][0] = 0;
        layer_1_weights[65][0] = 0;
        layer_1_weights[66][0] = 1;
        layer_1_weights[67][0] = 5;
        layer_1_weights[68][0] = 2;
        layer_1_weights[69][0] = 4;
        layer_1_weights[70][0] = 5;
        layer_1_weights[71][0] = 4;
        layer_1_weights[72][0] = 4;
        layer_1_weights[73][0] = 0;
        layer_1_weights[74][0] = 1;
        layer_1_weights[75][0] = 0;
        layer_1_weights[76][0] = 1;
        layer_1_weights[77][0] = 0;
        layer_1_weights[78][0] = -1;
        layer_1_weights[79][0] = 0;
        layer_1_weights[80][0] = 2;
        layer_1_weights[81][0] = 1;
        layer_1_weights[82][0] = 0;
        layer_1_weights[83][0] = 0;
        layer_1_weights[84][0] = -1;
        layer_1_weights[85][0] = 0;
        layer_1_weights[86][0] = 3;
        layer_1_weights[87][0] = 4;
        layer_1_weights[88][0] = 2;
        layer_1_weights[89][0] = 1;
        layer_1_weights[90][0] = 1;
        layer_1_weights[91][0] = 0;
        layer_1_weights[92][0] = -1;
        layer_1_weights[93][0] = 1;
        layer_1_weights[94][0] = -1;
        layer_1_weights[95][0] = -4;
        layer_1_weights[96][0] = 0;
        layer_1_weights[97][0] = 2;
        layer_1_weights[98][0] = 2;
        layer_1_weights[99][0] = 0;
        layer_1_weights[100][0] = 2;
        layer_1_weights[101][0] = 0;
        layer_1_weights[102][0] = 0;
        layer_1_weights[103][0] = 0;
        layer_1_weights[104][0] = 0;
        layer_1_weights[105][0] = -2;
        layer_1_weights[106][0] = -1;
        layer_1_weights[107][0] = 1;
        layer_1_weights[108][0] = 0;
        layer_1_weights[109][0] = 1;
        layer_1_weights[110][0] = -1;
        layer_1_weights[111][0] = 0;
        layer_1_weights[112][0] = 0;
        layer_1_weights[113][0] = 0;
        layer_1_weights[114][0] = 2;
        layer_1_weights[115][0] = 2;
        layer_1_weights[116][0] = 4;
        layer_1_weights[117][0] = 2;
        layer_1_weights[118][0] = 0;
        layer_1_weights[119][0] = -3;
        layer_1_weights[120][0] = 1;
        layer_1_weights[121][0] = 1;
        layer_1_weights[122][0] = 2;
        layer_1_weights[123][0] = 0;
        layer_1_weights[124][0] = -1;
        layer_1_weights[125][0] = -1;
        layer_1_weights[126][0] = 0;
        layer_1_weights[127][0] = 0;
        layer_1_weights[128][0] = -2;
        layer_1_weights[129][0] = -3;
        layer_1_weights[130][0] = -2;
        layer_1_weights[131][0] = -2;
        layer_1_weights[132][0] = -1;
        layer_1_weights[133][0] = -1;
        layer_1_weights[134][0] = -2;
        layer_1_weights[135][0] = -1;
        layer_1_weights[136][0] = -3;
        layer_1_weights[137][0] = -2;
        layer_1_weights[138][0] = 0;
        layer_1_weights[139][0] = 0;
        layer_1_weights[140][0] = 0;
        layer_1_weights[141][0] = 0;
        layer_1_weights[142][0] = 4;
        layer_1_weights[143][0] = -3;
        layer_1_weights[144][0] = 5;
        layer_1_weights[145][0] = 0;
        layer_1_weights[146][0] = 2;
        layer_1_weights[147][0] = 3;
        layer_1_weights[148][0] = -2;
        layer_1_weights[149][0] = -1;
        layer_1_weights[150][0] = 0;
        layer_1_weights[151][0] = 0;
        layer_1_weights[152][0] = 0;
        layer_1_weights[153][0] = 1;
        layer_1_weights[154][0] = 0;
        layer_1_weights[155][0] = 0;
        layer_1_weights[156][0] = -1;
        layer_1_weights[157][0] = -3;
        layer_1_weights[158][0] = -4;
        layer_1_weights[159][0] = -2;
        layer_1_weights[160][0] = -2;
        layer_1_weights[161][0] = -1;
        layer_1_weights[162][0] = -2;
        layer_1_weights[163][0] = -1;
        layer_1_weights[164][0] = -2;
        layer_1_weights[165][0] = -1;
        layer_1_weights[166][0] = 0;
        layer_1_weights[167][0] = 0;
        layer_1_weights[168][0] = 0;
        layer_1_weights[169][0] = 0;
        layer_1_weights[170][0] = -2;
        layer_1_weights[171][0] = -2;
        layer_1_weights[172][0] = 2;
        layer_1_weights[173][0] = 1;
        layer_1_weights[174][0] = 0;
        layer_1_weights[175][0] = 1;
        layer_1_weights[176][0] = -1;
        layer_1_weights[177][0] = -1;
        layer_1_weights[178][0] = -1;
        layer_1_weights[179][0] = 0;
        layer_1_weights[180][0] = 0;
        layer_1_weights[181][0] = -1;
        layer_1_weights[182][0] = -1;
        layer_1_weights[183][0] = 0;
        layer_1_weights[184][0] = -1;
        layer_1_weights[185][0] = -3;
        layer_1_weights[186][0] = -2;
        layer_1_weights[187][0] = -2;
        layer_1_weights[188][0] = -1;
        layer_1_weights[189][0] = 0;
        layer_1_weights[190][0] = -2;
        layer_1_weights[191][0] = -3;
        layer_1_weights[192][0] = -1;
        layer_1_weights[193][0] = -1;
        layer_1_weights[194][0] = -1;
        layer_1_weights[195][0] = -2;
        layer_1_weights[196][0] = 1;
        layer_1_weights[197][0] = 3;
        layer_1_weights[198][0] = -1;
        layer_1_weights[199][0] = 1;
        layer_1_weights[200][0] = 4;
        layer_1_weights[201][0] = 0;
        layer_1_weights[202][0] = 0;
        layer_1_weights[203][0] = 2;
        layer_1_weights[204][0] = -2;
        layer_1_weights[205][0] = 2;
        layer_1_weights[206][0] = 0;
        layer_1_weights[207][0] = -1;
        layer_1_weights[208][0] = 1;
        layer_1_weights[209][0] = -1;
        layer_1_weights[210][0] = 0;
        layer_1_weights[211][0] = -1;
        layer_1_weights[212][0] = -2;
        layer_1_weights[213][0] = -1;
        layer_1_weights[214][0] = -2;
        layer_1_weights[215][0] = -3;
        layer_1_weights[216][0] = -2;
        layer_1_weights[217][0] = 0;
        layer_1_weights[218][0] = -2;
        layer_1_weights[219][0] = -2;
        layer_1_weights[220][0] = -3;
        layer_1_weights[221][0] = -2;
        layer_1_weights[222][0] = -2;
        layer_1_weights[223][0] = -3;
        layer_1_weights[224][0] = 0;
        layer_1_weights[225][0] = 3;
        layer_1_weights[226][0] = 4;
        layer_1_weights[227][0] = 3;
        layer_1_weights[228][0] = 4;
        layer_1_weights[229][0] = 0;
        layer_1_weights[230][0] = 1;
        layer_1_weights[231][0] = 2;
        layer_1_weights[232][0] = 2;
        layer_1_weights[233][0] = 1;
        layer_1_weights[234][0] = -2;
        layer_1_weights[235][0] = 0;
        layer_1_weights[236][0] = -1;
        layer_1_weights[237][0] = 1;
        layer_1_weights[238][0] = -1;
        layer_1_weights[239][0] = 0;
        layer_1_weights[240][0] = -2;
        layer_1_weights[241][0] = -2;
        layer_1_weights[242][0] = -3;
        layer_1_weights[243][0] = -2;
        layer_1_weights[244][0] = 1;
        layer_1_weights[245][0] = 0;
        layer_1_weights[246][0] = -1;
        layer_1_weights[247][0] = -1;
        layer_1_weights[248][0] = -4;
        layer_1_weights[249][0] = -3;
        layer_1_weights[250][0] = -1;
        layer_1_weights[251][0] = -4;
        layer_1_weights[252][0] = 1;
        layer_1_weights[253][0] = 1;
        layer_1_weights[254][0] = 3;
        layer_1_weights[255][0] = 3;
        layer_1_weights[256][0] = 2;
        layer_1_weights[257][0] = 0;
        layer_1_weights[258][0] = 2;
        layer_1_weights[259][0] = 2;
        layer_1_weights[260][0] = 1;
        layer_1_weights[261][0] = 0;
        layer_1_weights[262][0] = 0;
        layer_1_weights[263][0] = 0;
        layer_1_weights[264][0] = 0;
        layer_1_weights[265][0] = 2;
        layer_1_weights[266][0] = 2;
        layer_1_weights[267][0] = -1;
        layer_1_weights[268][0] = -2;
        layer_1_weights[269][0] = -2;
        layer_1_weights[270][0] = -1;
        layer_1_weights[271][0] = -2;
        layer_1_weights[272][0] = 1;
        layer_1_weights[273][0] = 1;
        layer_1_weights[274][0] = -1;
        layer_1_weights[275][0] = -1;
        layer_1_weights[276][0] = 0;
        layer_1_weights[277][0] = -2;
        layer_1_weights[278][0] = -3;
        layer_1_weights[279][0] = 2;
        layer_1_weights[280][0] = 2;
        layer_1_weights[281][0] = 5;
        layer_1_weights[282][0] = -2;
        layer_1_weights[283][0] = -2;
        layer_1_weights[284][0] = 1;
        layer_1_weights[285][0] = 0;
        layer_1_weights[286][0] = -1;
        layer_1_weights[287][0] = 1;
        layer_1_weights[288][0] = 0;
        layer_1_weights[289][0] = 0;
        layer_1_weights[290][0] = 0;
        layer_1_weights[291][0] = 0;
        layer_1_weights[292][0] = 2;
        layer_1_weights[293][0] = 2;
        layer_1_weights[294][0] = 2;
        layer_1_weights[295][0] = 1;
        layer_1_weights[296][0] = 0;
        layer_1_weights[297][0] = -1;
        layer_1_weights[298][0] = -1;
        layer_1_weights[299][0] = -1;
        layer_1_weights[300][0] = -1;
        layer_1_weights[301][0] = 0;
        layer_1_weights[302][0] = 0;
        layer_1_weights[303][0] = 0;
        layer_1_weights[304][0] = 0;
        layer_1_weights[305][0] = -1;
        layer_1_weights[306][0] = -1;
        layer_1_weights[307][0] = 2;
        layer_1_weights[308][0] = 1;
        layer_1_weights[309][0] = 5;
        layer_1_weights[310][0] = -1;
        layer_1_weights[311][0] = 0;
        layer_1_weights[312][0] = 1;
        layer_1_weights[313][0] = -1;
        layer_1_weights[314][0] = -2;
        layer_1_weights[315][0] = 1;
        layer_1_weights[316][0] = -1;
        layer_1_weights[317][0] = 0;
        layer_1_weights[318][0] = 0;
        layer_1_weights[319][0] = -1;
        layer_1_weights[320][0] = 1;
        layer_1_weights[321][0] = 1;
        layer_1_weights[322][0] = 1;
        layer_1_weights[323][0] = 0;
        layer_1_weights[324][0] = -1;
        layer_1_weights[325][0] = 1;
        layer_1_weights[326][0] = -1;
        layer_1_weights[327][0] = 0;
        layer_1_weights[328][0] = 0;
        layer_1_weights[329][0] = 0;
        layer_1_weights[330][0] = 1;
        layer_1_weights[331][0] = 2;
        layer_1_weights[332][0] = -2;
        layer_1_weights[333][0] = -3;
        layer_1_weights[334][0] = -1;
        layer_1_weights[335][0] = -2;
        layer_1_weights[336][0] = 1;
        layer_1_weights[337][0] = 5;
        layer_1_weights[338][0] = -1;
        layer_1_weights[339][0] = 1;
        layer_1_weights[340][0] = 2;
        layer_1_weights[341][0] = 1;
        layer_1_weights[342][0] = 0;
        layer_1_weights[343][0] = 1;
        layer_1_weights[344][0] = 2;
        layer_1_weights[345][0] = 0;
        layer_1_weights[346][0] = 0;
        layer_1_weights[347][0] = -1;
        layer_1_weights[348][0] = 0;
        layer_1_weights[349][0] = 0;
        layer_1_weights[350][0] = 0;
        layer_1_weights[351][0] = 1;
        layer_1_weights[352][0] = 2;
        layer_1_weights[353][0] = 0;
        layer_1_weights[354][0] = 0;
        layer_1_weights[355][0] = 0;
        layer_1_weights[356][0] = 0;
        layer_1_weights[357][0] = 0;
        layer_1_weights[358][0] = 2;
        layer_1_weights[359][0] = 1;
        layer_1_weights[360][0] = 1;
        layer_1_weights[361][0] = -2;
        layer_1_weights[362][0] = -5;
        layer_1_weights[363][0] = -3;
        layer_1_weights[364][0] = 0;
        layer_1_weights[365][0] = 3;
        layer_1_weights[366][0] = 1;
        layer_1_weights[367][0] = 2;
        layer_1_weights[368][0] = 0;
        layer_1_weights[369][0] = 1;
        layer_1_weights[370][0] = 2;
        layer_1_weights[371][0] = -1;
        layer_1_weights[372][0] = -1;
        layer_1_weights[373][0] = 1;
        layer_1_weights[374][0] = 0;
        layer_1_weights[375][0] = 0;
        layer_1_weights[376][0] = -1;
        layer_1_weights[377][0] = -1;
        layer_1_weights[378][0] = 0;
        layer_1_weights[379][0] = 4;
        layer_1_weights[380][0] = 2;
        layer_1_weights[381][0] = 1;
        layer_1_weights[382][0] = 0;
        layer_1_weights[383][0] = 0;
        layer_1_weights[384][0] = 0;
        layer_1_weights[385][0] = 1;
        layer_1_weights[386][0] = 3;
        layer_1_weights[387][0] = 0;
        layer_1_weights[388][0] = 3;
        layer_1_weights[389][0] = -2;
        layer_1_weights[390][0] = -4;
        layer_1_weights[391][0] = 0;
        layer_1_weights[392][0] = -1;
        layer_1_weights[393][0] = 2;
        layer_1_weights[394][0] = 4;
        layer_1_weights[395][0] = 5;
        layer_1_weights[396][0] = -1;
        layer_1_weights[397][0] = 1;
        layer_1_weights[398][0] = 0;
        layer_1_weights[399][0] = -1;
        layer_1_weights[400][0] = 0;
        layer_1_weights[401][0] = 0;
        layer_1_weights[402][0] = -1;
        layer_1_weights[403][0] = -1;
        layer_1_weights[404][0] = -1;
        layer_1_weights[405][0] = -2;
        layer_1_weights[406][0] = 1;
        layer_1_weights[407][0] = 2;
        layer_1_weights[408][0] = 1;
        layer_1_weights[409][0] = 0;
        layer_1_weights[410][0] = -1;
        layer_1_weights[411][0] = 1;
        layer_1_weights[412][0] = 1;
        layer_1_weights[413][0] = 1;
        layer_1_weights[414][0] = 4;
        layer_1_weights[415][0] = 3;
        layer_1_weights[416][0] = 1;
        layer_1_weights[417][0] = 1;
        layer_1_weights[418][0] = -3;
        layer_1_weights[419][0] = 1;
        layer_1_weights[420][0] = -1;
        layer_1_weights[421][0] = 0;
        layer_1_weights[422][0] = 3;
        layer_1_weights[423][0] = 4;
        layer_1_weights[424][0] = -1;
        layer_1_weights[425][0] = -1;
        layer_1_weights[426][0] = 1;
        layer_1_weights[427][0] = 0;
        layer_1_weights[428][0] = 0;
        layer_1_weights[429][0] = -1;
        layer_1_weights[430][0] = -1;
        layer_1_weights[431][0] = -3;
        layer_1_weights[432][0] = -4;
        layer_1_weights[433][0] = 1;
        layer_1_weights[434][0] = 4;
        layer_1_weights[435][0] = 1;
        layer_1_weights[436][0] = 2;
        layer_1_weights[437][0] = -1;
        layer_1_weights[438][0] = -1;
        layer_1_weights[439][0] = 1;
        layer_1_weights[440][0] = 0;
        layer_1_weights[441][0] = 0;
        layer_1_weights[442][0] = 2;
        layer_1_weights[443][0] = 1;
        layer_1_weights[444][0] = -1;
        layer_1_weights[445][0] = 2;
        layer_1_weights[446][0] = -3;
        layer_1_weights[447][0] = -2;
        layer_1_weights[448][0] = 2;
        layer_1_weights[449][0] = 0;
        layer_1_weights[450][0] = 3;
        layer_1_weights[451][0] = 2;
        layer_1_weights[452][0] = -3;
        layer_1_weights[453][0] = 1;
        layer_1_weights[454][0] = 1;
        layer_1_weights[455][0] = 0;
        layer_1_weights[456][0] = -2;
        layer_1_weights[457][0] = 0;
        layer_1_weights[458][0] = -1;
        layer_1_weights[459][0] = -3;
        layer_1_weights[460][0] = -3;
        layer_1_weights[461][0] = 3;
        layer_1_weights[462][0] = 4;
        layer_1_weights[463][0] = 2;
        layer_1_weights[464][0] = 1;
        layer_1_weights[465][0] = 0;
        layer_1_weights[466][0] = -1;
        layer_1_weights[467][0] = 0;
        layer_1_weights[468][0] = 0;
        layer_1_weights[469][0] = 0;
        layer_1_weights[470][0] = 1;
        layer_1_weights[471][0] = 0;
        layer_1_weights[472][0] = 1;
        layer_1_weights[473][0] = 2;
        layer_1_weights[474][0] = -4;
        layer_1_weights[475][0] = -3;
        layer_1_weights[476][0] = 0;
        layer_1_weights[477][0] = 1;
        layer_1_weights[478][0] = 0;
        layer_1_weights[479][0] = 2;
        layer_1_weights[480][0] = 0;
        layer_1_weights[481][0] = 0;
        layer_1_weights[482][0] = 0;
        layer_1_weights[483][0] = 0;
        layer_1_weights[484][0] = -1;
        layer_1_weights[485][0] = -2;
        layer_1_weights[486][0] = -2;
        layer_1_weights[487][0] = -3;
        layer_1_weights[488][0] = -1;
        layer_1_weights[489][0] = 3;
        layer_1_weights[490][0] = 5;
        layer_1_weights[491][0] = 3;
        layer_1_weights[492][0] = 1;
        layer_1_weights[493][0] = 0;
        layer_1_weights[494][0] = 1;
        layer_1_weights[495][0] = 1;
        layer_1_weights[496][0] = 0;
        layer_1_weights[497][0] = 0;
        layer_1_weights[498][0] = 1;
        layer_1_weights[499][0] = -1;
        layer_1_weights[500][0] = 2;
        layer_1_weights[501][0] = 2;
        layer_1_weights[502][0] = 0;
        layer_1_weights[503][0] = -1;
        layer_1_weights[504][0] = 1;
        layer_1_weights[505][0] = 1;
        layer_1_weights[506][0] = 4;
        layer_1_weights[507][0] = -2;
        layer_1_weights[508][0] = 0;
        layer_1_weights[509][0] = 0;
        layer_1_weights[510][0] = -1;
        layer_1_weights[511][0] = 0;
        layer_1_weights[512][0] = -3;
        layer_1_weights[513][0] = -4;
        layer_1_weights[514][0] = -4;
        layer_1_weights[515][0] = -1;
        layer_1_weights[516][0] = 1;
        layer_1_weights[517][0] = 3;
        layer_1_weights[518][0] = 4;
        layer_1_weights[519][0] = 1;
        layer_1_weights[520][0] = 0;
        layer_1_weights[521][0] = 1;
        layer_1_weights[522][0] = 3;
        layer_1_weights[523][0] = 1;
        layer_1_weights[524][0] = 3;
        layer_1_weights[525][0] = -1;
        layer_1_weights[526][0] = 2;
        layer_1_weights[527][0] = 0;
        layer_1_weights[528][0] = 1;
        layer_1_weights[529][0] = 2;
        layer_1_weights[530][0] = 4;
        layer_1_weights[531][0] = 3;
        layer_1_weights[532][0] = 0;
        layer_1_weights[533][0] = 3;
        layer_1_weights[534][0] = 2;
        layer_1_weights[535][0] = -2;
        layer_1_weights[536][0] = -4;
        layer_1_weights[537][0] = -3;
        layer_1_weights[538][0] = -1;
        layer_1_weights[539][0] = -2;
        layer_1_weights[540][0] = -3;
        layer_1_weights[541][0] = -2;
        layer_1_weights[542][0] = -2;
        layer_1_weights[543][0] = -2;
        layer_1_weights[544][0] = 2;
        layer_1_weights[545][0] = 4;
        layer_1_weights[546][0] = 3;
        layer_1_weights[547][0] = 2;
        layer_1_weights[548][0] = 1;
        layer_1_weights[549][0] = 1;
        layer_1_weights[550][0] = 1;
        layer_1_weights[551][0] = 2;
        layer_1_weights[552][0] = 1;
        layer_1_weights[553][0] = 0;
        layer_1_weights[554][0] = -1;
        layer_1_weights[555][0] = 0;
        layer_1_weights[556][0] = 3;
        layer_1_weights[557][0] = 1;
        layer_1_weights[558][0] = 0;
        layer_1_weights[559][0] = 2;
        layer_1_weights[560][0] = 0;
        layer_1_weights[561][0] = 1;
        layer_1_weights[562][0] = -1;
        layer_1_weights[563][0] = 0;
        layer_1_weights[564][0] = -2;
        layer_1_weights[565][0] = -4;
        layer_1_weights[566][0] = 0;
        layer_1_weights[567][0] = -1;
        layer_1_weights[568][0] = -4;
        layer_1_weights[569][0] = -2;
        layer_1_weights[570][0] = -1;
        layer_1_weights[571][0] = 1;
        layer_1_weights[572][0] = 3;
        layer_1_weights[573][0] = 3;
        layer_1_weights[574][0] = 2;
        layer_1_weights[575][0] = 2;
        layer_1_weights[576][0] = 1;
        layer_1_weights[577][0] = 1;
        layer_1_weights[578][0] = 3;
        layer_1_weights[579][0] = 1;
        layer_1_weights[580][0] = 1;
        layer_1_weights[581][0] = -2;
        layer_1_weights[582][0] = -3;
        layer_1_weights[583][0] = -2;
        layer_1_weights[584][0] = 0;
        layer_1_weights[585][0] = -1;
        layer_1_weights[586][0] = 2;
        layer_1_weights[587][0] = 1;
        layer_1_weights[588][0] = 0;
        layer_1_weights[589][0] = -2;
        layer_1_weights[590][0] = -2;
        layer_1_weights[591][0] = -1;
        layer_1_weights[592][0] = 0;
        layer_1_weights[593][0] = 1;
        layer_1_weights[594][0] = 0;
        layer_1_weights[595][0] = 1;
        layer_1_weights[596][0] = -1;
        layer_1_weights[597][0] = -1;
        layer_1_weights[598][0] = -1;
        layer_1_weights[599][0] = 0;
        layer_1_weights[600][0] = 1;
        layer_1_weights[601][0] = 2;
        layer_1_weights[602][0] = 2;
        layer_1_weights[603][0] = 3;
        layer_1_weights[604][0] = 1;
        layer_1_weights[605][0] = 2;
        layer_1_weights[606][0] = 2;
        layer_1_weights[607][0] = 0;
        layer_1_weights[608][0] = 0;
        layer_1_weights[609][0] = 1;
        layer_1_weights[610][0] = -4;
        layer_1_weights[611][0] = -1;
        layer_1_weights[612][0] = -1;
        layer_1_weights[613][0] = 1;
        layer_1_weights[614][0] = 4;
        layer_1_weights[615][0] = 0;
        layer_1_weights[616][0] = 1;
        layer_1_weights[617][0] = 0;
        layer_1_weights[618][0] = -1;
        layer_1_weights[619][0] = -1;
        layer_1_weights[620][0] = 2;
        layer_1_weights[621][0] = 1;
        layer_1_weights[622][0] = -1;
        layer_1_weights[623][0] = 0;
        layer_1_weights[624][0] = 1;
        layer_1_weights[625][0] = 1;
        layer_1_weights[626][0] = -1;
        layer_1_weights[627][0] = -3;
        layer_1_weights[628][0] = -1;
        layer_1_weights[629][0] = -1;
        layer_1_weights[630][0] = 1;
        layer_1_weights[631][0] = 2;
        layer_1_weights[632][0] = 1;
        layer_1_weights[633][0] = 1;
        layer_1_weights[634][0] = 0;
        layer_1_weights[635][0] = -1;
        layer_1_weights[636][0] = 0;
        layer_1_weights[637][0] = 0;
        layer_1_weights[638][0] = 0;
        layer_1_weights[639][0] = -7;
        layer_1_weights[640][0] = -1;
        layer_1_weights[641][0] = 2;
        layer_1_weights[642][0] = 2;
        layer_1_weights[643][0] = 0;
        layer_1_weights[644][0] = 0;
        layer_1_weights[645][0] = 0;
        layer_1_weights[646][0] = -2;
        layer_1_weights[647][0] = -3;
        layer_1_weights[648][0] = -5;
        layer_1_weights[649][0] = -1;
        layer_1_weights[650][0] = -1;
        layer_1_weights[651][0] = -3;
        layer_1_weights[652][0] = -4;
        layer_1_weights[653][0] = -1;
        layer_1_weights[654][0] = -3;
        layer_1_weights[655][0] = -3;
        layer_1_weights[656][0] = -1;
        layer_1_weights[657][0] = -1;
        layer_1_weights[658][0] = 0;
        layer_1_weights[659][0] = -1;
        layer_1_weights[660][0] = 1;
        layer_1_weights[661][0] = 0;
        layer_1_weights[662][0] = 1;
        layer_1_weights[663][0] = 0;
        layer_1_weights[664][0] = 0;
        layer_1_weights[665][0] = -1;
        layer_1_weights[666][0] = -3;
        layer_1_weights[667][0] = -9;
        layer_1_weights[668][0] = -6;
        layer_1_weights[669][0] = -4;
        layer_1_weights[670][0] = 3;
        layer_1_weights[671][0] = 0;
        layer_1_weights[672][0] = 0;
        layer_1_weights[673][0] = 1;
        layer_1_weights[674][0] = 1;
        layer_1_weights[675][0] = 2;
        layer_1_weights[676][0] = -2;
        layer_1_weights[677][0] = 0;
        layer_1_weights[678][0] = 0;
        layer_1_weights[679][0] = 2;
        layer_1_weights[680][0] = 0;
        layer_1_weights[681][0] = 0;
        layer_1_weights[682][0] = -2;
        layer_1_weights[683][0] = -1;
        layer_1_weights[684][0] = -2;
        layer_1_weights[685][0] = -1;
        layer_1_weights[686][0] = -1;
        layer_1_weights[687][0] = 1;
        layer_1_weights[688][0] = -1;
        layer_1_weights[689][0] = -1;
        layer_1_weights[690][0] = -1;
        layer_1_weights[691][0] = -3;
        layer_1_weights[692][0] = -2;
        layer_1_weights[693][0] = -2;
        layer_1_weights[694][0] = -3;
        layer_1_weights[695][0] = -9;
        layer_1_weights[696][0] = -4;
        layer_1_weights[697][0] = 1;
        layer_1_weights[698][0] = 0;
        layer_1_weights[699][0] = 0;
        layer_1_weights[700][0] = 0;
        layer_1_weights[701][0] = 0;
        layer_1_weights[702][0] = -2;
        layer_1_weights[703][0] = 1;
        layer_1_weights[704][0] = -2;
        layer_1_weights[705][0] = -2;
        layer_1_weights[706][0] = -1;
        layer_1_weights[707][0] = 1;
        layer_1_weights[708][0] = 2;
        layer_1_weights[709][0] = -1;
        layer_1_weights[710][0] = -4;
        layer_1_weights[711][0] = -2;
        layer_1_weights[712][0] = -2;
        layer_1_weights[713][0] = -3;
        layer_1_weights[714][0] = -3;
        layer_1_weights[715][0] = -2;
        layer_1_weights[716][0] = -2;
        layer_1_weights[717][0] = -2;
        layer_1_weights[718][0] = -4;
        layer_1_weights[719][0] = -3;
        layer_1_weights[720][0] = -4;
        layer_1_weights[721][0] = -2;
        layer_1_weights[722][0] = -1;
        layer_1_weights[723][0] = 0;
        layer_1_weights[724][0] = -1;
        layer_1_weights[725][0] = -2;
        layer_1_weights[726][0] = 0;
        layer_1_weights[727][0] = 0;
        layer_1_weights[728][0] = 0;
        layer_1_weights[729][0] = 0;
        layer_1_weights[730][0] = 1;
        layer_1_weights[731][0] = -2;
        layer_1_weights[732][0] = -3;
        layer_1_weights[733][0] = -1;
        layer_1_weights[734][0] = -1;
        layer_1_weights[735][0] = 0;
        layer_1_weights[736][0] = 0;
        layer_1_weights[737][0] = -1;
        layer_1_weights[738][0] = -2;
        layer_1_weights[739][0] = -3;
        layer_1_weights[740][0] = -2;
        layer_1_weights[741][0] = -2;
        layer_1_weights[742][0] = -3;
        layer_1_weights[743][0] = -3;
        layer_1_weights[744][0] = -1;
        layer_1_weights[745][0] = -1;
        layer_1_weights[746][0] = -2;
        layer_1_weights[747][0] = -2;
        layer_1_weights[748][0] = -1;
        layer_1_weights[749][0] = 0;
        layer_1_weights[750][0] = -2;
        layer_1_weights[751][0] = -1;
        layer_1_weights[752][0] = 1;
        layer_1_weights[753][0] = 2;
        layer_1_weights[754][0] = 1;
        layer_1_weights[755][0] = 0;
        layer_1_weights[756][0] = 0;
        layer_1_weights[757][0] = 0;
        layer_1_weights[758][0] = 0;
        layer_1_weights[759][0] = 0;
        layer_1_weights[760][0] = 2;
        layer_1_weights[761][0] = 4;
        layer_1_weights[762][0] = 2;
        layer_1_weights[763][0] = 4;
        layer_1_weights[764][0] = 4;
        layer_1_weights[765][0] = 1;
        layer_1_weights[766][0] = 0;
        layer_1_weights[767][0] = -1;
        layer_1_weights[768][0] = 0;
        layer_1_weights[769][0] = 1;
        layer_1_weights[770][0] = -4;
        layer_1_weights[771][0] = -3;
        layer_1_weights[772][0] = 0;
        layer_1_weights[773][0] = 3;
        layer_1_weights[774][0] = 3;
        layer_1_weights[775][0] = 3;
        layer_1_weights[776][0] = 0;
        layer_1_weights[777][0] = 2;
        layer_1_weights[778][0] = 1;
        layer_1_weights[779][0] = 2;
        layer_1_weights[780][0] = 0;
        layer_1_weights[781][0] = 0;
        layer_1_weights[782][0] = 0;
        layer_1_weights[783][0] = -1;
        layer_1_weights[0][1] = 0;
        layer_1_weights[1][1] = 0;
        layer_1_weights[2][1] = 0;
        layer_1_weights[3][1] = 0;
        layer_1_weights[4][1] = 0;
        layer_1_weights[5][1] = 1;
        layer_1_weights[6][1] = 0;
        layer_1_weights[7][1] = -1;
        layer_1_weights[8][1] = 0;
        layer_1_weights[9][1] = 0;
        layer_1_weights[10][1] = 0;
        layer_1_weights[11][1] = 0;
        layer_1_weights[12][1] = 1;
        layer_1_weights[13][1] = 1;
        layer_1_weights[14][1] = 0;
        layer_1_weights[15][1] = 0;
        layer_1_weights[16][1] = 0;
        layer_1_weights[17][1] = 0;
        layer_1_weights[18][1] = 0;
        layer_1_weights[19][1] = 0;
        layer_1_weights[20][1] = 0;
        layer_1_weights[21][1] = 0;
        layer_1_weights[22][1] = 0;
        layer_1_weights[23][1] = 0;
        layer_1_weights[24][1] = -1;
        layer_1_weights[25][1] = -1;
        layer_1_weights[26][1] = 0;
        layer_1_weights[27][1] = 0;
        layer_1_weights[28][1] = -1;
        layer_1_weights[29][1] = 1;
        layer_1_weights[30][1] = 0;
        layer_1_weights[31][1] = 0;
        layer_1_weights[32][1] = -1;
        layer_1_weights[33][1] = 0;
        layer_1_weights[34][1] = 0;
        layer_1_weights[35][1] = 0;
        layer_1_weights[36][1] = 0;
        layer_1_weights[37][1] = -1;
        layer_1_weights[38][1] = -1;
        layer_1_weights[39][1] = 3;
        layer_1_weights[40][1] = 0;
        layer_1_weights[41][1] = 2;
        layer_1_weights[42][1] = -3;
        layer_1_weights[43][1] = 2;
        layer_1_weights[44][1] = 1;
        layer_1_weights[45][1] = 2;
        layer_1_weights[46][1] = -2;
        layer_1_weights[47][1] = 1;
        layer_1_weights[48][1] = 2;
        layer_1_weights[49][1] = 0;
        layer_1_weights[50][1] = 2;
        layer_1_weights[51][1] = 1;
        layer_1_weights[52][1] = 0;
        layer_1_weights[53][1] = 0;
        layer_1_weights[54][1] = 0;
        layer_1_weights[55][1] = 0;
        layer_1_weights[56][1] = 0;
        layer_1_weights[57][1] = -1;
        layer_1_weights[58][1] = 0;
        layer_1_weights[59][1] = 0;
        layer_1_weights[60][1] = 0;
        layer_1_weights[61][1] = -2;
        layer_1_weights[62][1] = 0;
        layer_1_weights[63][1] = -1;
        layer_1_weights[64][1] = 3;
        layer_1_weights[65][1] = 3;
        layer_1_weights[66][1] = 2;
        layer_1_weights[67][1] = 0;
        layer_1_weights[68][1] = -2;
        layer_1_weights[69][1] = -4;
        layer_1_weights[70][1] = -6;
        layer_1_weights[71][1] = -4;
        layer_1_weights[72][1] = -3;
        layer_1_weights[73][1] = 0;
        layer_1_weights[74][1] = 1;
        layer_1_weights[75][1] = 1;
        layer_1_weights[76][1] = -1;
        layer_1_weights[77][1] = 1;
        layer_1_weights[78][1] = 0;
        layer_1_weights[79][1] = 2;
        layer_1_weights[80][1] = -2;
        layer_1_weights[81][1] = 0;
        layer_1_weights[82][1] = 0;
        layer_1_weights[83][1] = 1;
        layer_1_weights[84][1] = -1;
        layer_1_weights[85][1] = 0;
        layer_1_weights[86][1] = 0;
        layer_1_weights[87][1] = 1;
        layer_1_weights[88][1] = 0;
        layer_1_weights[89][1] = 2;
        layer_1_weights[90][1] = -1;
        layer_1_weights[91][1] = 0;
        layer_1_weights[92][1] = 4;
        layer_1_weights[93][1] = 1;
        layer_1_weights[94][1] = 1;
        layer_1_weights[95][1] = 3;
        layer_1_weights[96][1] = 1;
        layer_1_weights[97][1] = 1;
        layer_1_weights[98][1] = 0;
        layer_1_weights[99][1] = 1;
        layer_1_weights[100][1] = -1;
        layer_1_weights[101][1] = -1;
        layer_1_weights[102][1] = -1;
        layer_1_weights[103][1] = -1;
        layer_1_weights[104][1] = 1;
        layer_1_weights[105][1] = 2;
        layer_1_weights[106][1] = 1;
        layer_1_weights[107][1] = -1;
        layer_1_weights[108][1] = 6;
        layer_1_weights[109][1] = 3;
        layer_1_weights[110][1] = 1;
        layer_1_weights[111][1] = 1;
        layer_1_weights[112][1] = 0;
        layer_1_weights[113][1] = 1;
        layer_1_weights[114][1] = 2;
        layer_1_weights[115][1] = 1;
        layer_1_weights[116][1] = -2;
        layer_1_weights[117][1] = 1;
        layer_1_weights[118][1] = 0;
        layer_1_weights[119][1] = 0;
        layer_1_weights[120][1] = -1;
        layer_1_weights[121][1] = -2;
        layer_1_weights[122][1] = 0;
        layer_1_weights[123][1] = 2;
        layer_1_weights[124][1] = 1;
        layer_1_weights[125][1] = 1;
        layer_1_weights[126][1] = -1;
        layer_1_weights[127][1] = 0;
        layer_1_weights[128][1] = 0;
        layer_1_weights[129][1] = -1;
        layer_1_weights[130][1] = -1;
        layer_1_weights[131][1] = 0;
        layer_1_weights[132][1] = -1;
        layer_1_weights[133][1] = -1;
        layer_1_weights[134][1] = 1;
        layer_1_weights[135][1] = -3;
        layer_1_weights[136][1] = 2;
        layer_1_weights[137][1] = 2;
        layer_1_weights[138][1] = 2;
        layer_1_weights[139][1] = -1;
        layer_1_weights[140][1] = -1;
        layer_1_weights[141][1] = 0;
        layer_1_weights[142][1] = -3;
        layer_1_weights[143][1] = 1;
        layer_1_weights[144][1] = -3;
        layer_1_weights[145][1] = -1;
        layer_1_weights[146][1] = 0;
        layer_1_weights[147][1] = 3;
        layer_1_weights[148][1] = 1;
        layer_1_weights[149][1] = 1;
        layer_1_weights[150][1] = 1;
        layer_1_weights[151][1] = 1;
        layer_1_weights[152][1] = 2;
        layer_1_weights[153][1] = 1;
        layer_1_weights[154][1] = 0;
        layer_1_weights[155][1] = 1;
        layer_1_weights[156][1] = -1;
        layer_1_weights[157][1] = -1;
        layer_1_weights[158][1] = -1;
        layer_1_weights[159][1] = -1;
        layer_1_weights[160][1] = 0;
        layer_1_weights[161][1] = -2;
        layer_1_weights[162][1] = -1;
        layer_1_weights[163][1] = -3;
        layer_1_weights[164][1] = -3;
        layer_1_weights[165][1] = 5;
        layer_1_weights[166][1] = 2;
        layer_1_weights[167][1] = 2;
        layer_1_weights[168][1] = 0;
        layer_1_weights[169][1] = 0;
        layer_1_weights[170][1] = 3;
        layer_1_weights[171][1] = 4;
        layer_1_weights[172][1] = 0;
        layer_1_weights[173][1] = 2;
        layer_1_weights[174][1] = 0;
        layer_1_weights[175][1] = 3;
        layer_1_weights[176][1] = 2;
        layer_1_weights[177][1] = 2;
        layer_1_weights[178][1] = 2;
        layer_1_weights[179][1] = 2;
        layer_1_weights[180][1] = 4;
        layer_1_weights[181][1] = 1;
        layer_1_weights[182][1] = 2;
        layer_1_weights[183][1] = 2;
        layer_1_weights[184][1] = 1;
        layer_1_weights[185][1] = 1;
        layer_1_weights[186][1] = -1;
        layer_1_weights[187][1] = 1;
        layer_1_weights[188][1] = 0;
        layer_1_weights[189][1] = 0;
        layer_1_weights[190][1] = -1;
        layer_1_weights[191][1] = -2;
        layer_1_weights[192][1] = -1;
        layer_1_weights[193][1] = 1;
        layer_1_weights[194][1] = 1;
        layer_1_weights[195][1] = 0;
        layer_1_weights[196][1] = 0;
        layer_1_weights[197][1] = 4;
        layer_1_weights[198][1] = 3;
        layer_1_weights[199][1] = 0;
        layer_1_weights[200][1] = -3;
        layer_1_weights[201][1] = -2;
        layer_1_weights[202][1] = 1;
        layer_1_weights[203][1] = 1;
        layer_1_weights[204][1] = 2;
        layer_1_weights[205][1] = 0;
        layer_1_weights[206][1] = 2;
        layer_1_weights[207][1] = 1;
        layer_1_weights[208][1] = 1;
        layer_1_weights[209][1] = 1;
        layer_1_weights[210][1] = 1;
        layer_1_weights[211][1] = 3;
        layer_1_weights[212][1] = 2;
        layer_1_weights[213][1] = 0;
        layer_1_weights[214][1] = 0;
        layer_1_weights[215][1] = 0;
        layer_1_weights[216][1] = 0;
        layer_1_weights[217][1] = 1;
        layer_1_weights[218][1] = 0;
        layer_1_weights[219][1] = 1;
        layer_1_weights[220][1] = -1;
        layer_1_weights[221][1] = -1;
        layer_1_weights[222][1] = -3;
        layer_1_weights[223][1] = 1;
        layer_1_weights[224][1] = -2;
        layer_1_weights[225][1] = 0;
        layer_1_weights[226][1] = -1;
        layer_1_weights[227][1] = 1;
        layer_1_weights[228][1] = 0;
        layer_1_weights[229][1] = 2;
        layer_1_weights[230][1] = 1;
        layer_1_weights[231][1] = 1;
        layer_1_weights[232][1] = 2;
        layer_1_weights[233][1] = 1;
        layer_1_weights[234][1] = 0;
        layer_1_weights[235][1] = 1;
        layer_1_weights[236][1] = 1;
        layer_1_weights[237][1] = 2;
        layer_1_weights[238][1] = 3;
        layer_1_weights[239][1] = 1;
        layer_1_weights[240][1] = 1;
        layer_1_weights[241][1] = 2;
        layer_1_weights[242][1] = 1;
        layer_1_weights[243][1] = 2;
        layer_1_weights[244][1] = 0;
        layer_1_weights[245][1] = 0;
        layer_1_weights[246][1] = -1;
        layer_1_weights[247][1] = -1;
        layer_1_weights[248][1] = 1;
        layer_1_weights[249][1] = 0;
        layer_1_weights[250][1] = -2;
        layer_1_weights[251][1] = 5;
        layer_1_weights[252][1] = 3;
        layer_1_weights[253][1] = 1;
        layer_1_weights[254][1] = 1;
        layer_1_weights[255][1] = 4;
        layer_1_weights[256][1] = 2;
        layer_1_weights[257][1] = 3;
        layer_1_weights[258][1] = 2;
        layer_1_weights[259][1] = 3;
        layer_1_weights[260][1] = 2;
        layer_1_weights[261][1] = 2;
        layer_1_weights[262][1] = 3;
        layer_1_weights[263][1] = 1;
        layer_1_weights[264][1] = 2;
        layer_1_weights[265][1] = 2;
        layer_1_weights[266][1] = 2;
        layer_1_weights[267][1] = 1;
        layer_1_weights[268][1] = 1;
        layer_1_weights[269][1] = 1;
        layer_1_weights[270][1] = 1;
        layer_1_weights[271][1] = 0;
        layer_1_weights[272][1] = 2;
        layer_1_weights[273][1] = 1;
        layer_1_weights[274][1] = 0;
        layer_1_weights[275][1] = -1;
        layer_1_weights[276][1] = 2;
        layer_1_weights[277][1] = 3;
        layer_1_weights[278][1] = 3;
        layer_1_weights[279][1] = 4;
        layer_1_weights[280][1] = 3;
        layer_1_weights[281][1] = 0;
        layer_1_weights[282][1] = 2;
        layer_1_weights[283][1] = 4;
        layer_1_weights[284][1] = 1;
        layer_1_weights[285][1] = 3;
        layer_1_weights[286][1] = 5;
        layer_1_weights[287][1] = 1;
        layer_1_weights[288][1] = 2;
        layer_1_weights[289][1] = 2;
        layer_1_weights[290][1] = 2;
        layer_1_weights[291][1] = 2;
        layer_1_weights[292][1] = 0;
        layer_1_weights[293][1] = 3;
        layer_1_weights[294][1] = 2;
        layer_1_weights[295][1] = 2;
        layer_1_weights[296][1] = -1;
        layer_1_weights[297][1] = 1;
        layer_1_weights[298][1] = 0;
        layer_1_weights[299][1] = 1;
        layer_1_weights[300][1] = 1;
        layer_1_weights[301][1] = 2;
        layer_1_weights[302][1] = 0;
        layer_1_weights[303][1] = -1;
        layer_1_weights[304][1] = 2;
        layer_1_weights[305][1] = 5;
        layer_1_weights[306][1] = 6;
        layer_1_weights[307][1] = 0;
        layer_1_weights[308][1] = 2;
        layer_1_weights[309][1] = 1;
        layer_1_weights[310][1] = 2;
        layer_1_weights[311][1] = 1;
        layer_1_weights[312][1] = 4;
        layer_1_weights[313][1] = 1;
        layer_1_weights[314][1] = 3;
        layer_1_weights[315][1] = 3;
        layer_1_weights[316][1] = 1;
        layer_1_weights[317][1] = 1;
        layer_1_weights[318][1] = 0;
        layer_1_weights[319][1] = 1;
        layer_1_weights[320][1] = 0;
        layer_1_weights[321][1] = 2;
        layer_1_weights[322][1] = 3;
        layer_1_weights[323][1] = 0;
        layer_1_weights[324][1] = 0;
        layer_1_weights[325][1] = 0;
        layer_1_weights[326][1] = 2;
        layer_1_weights[327][1] = 2;
        layer_1_weights[328][1] = 2;
        layer_1_weights[329][1] = 0;
        layer_1_weights[330][1] = -1;
        layer_1_weights[331][1] = 0;
        layer_1_weights[332][1] = 1;
        layer_1_weights[333][1] = 3;
        layer_1_weights[334][1] = 4;
        layer_1_weights[335][1] = 1;
        layer_1_weights[336][1] = 0;
        layer_1_weights[337][1] = 4;
        layer_1_weights[338][1] = 2;
        layer_1_weights[339][1] = 2;
        layer_1_weights[340][1] = 4;
        layer_1_weights[341][1] = 3;
        layer_1_weights[342][1] = 3;
        layer_1_weights[343][1] = 1;
        layer_1_weights[344][1] = 1;
        layer_1_weights[345][1] = -1;
        layer_1_weights[346][1] = 0;
        layer_1_weights[347][1] = 0;
        layer_1_weights[348][1] = -1;
        layer_1_weights[349][1] = 0;
        layer_1_weights[350][1] = 1;
        layer_1_weights[351][1] = 1;
        layer_1_weights[352][1] = 1;
        layer_1_weights[353][1] = 1;
        layer_1_weights[354][1] = 1;
        layer_1_weights[355][1] = 1;
        layer_1_weights[356][1] = 1;
        layer_1_weights[357][1] = -2;
        layer_1_weights[358][1] = -3;
        layer_1_weights[359][1] = 0;
        layer_1_weights[360][1] = -3;
        layer_1_weights[361][1] = -2;
        layer_1_weights[362][1] = -1;
        layer_1_weights[363][1] = 1;
        layer_1_weights[364][1] = 1;
        layer_1_weights[365][1] = 1;
        layer_1_weights[366][1] = -1;
        layer_1_weights[367][1] = 1;
        layer_1_weights[368][1] = 3;
        layer_1_weights[369][1] = 1;
        layer_1_weights[370][1] = -2;
        layer_1_weights[371][1] = -1;
        layer_1_weights[372][1] = -1;
        layer_1_weights[373][1] = -2;
        layer_1_weights[374][1] = -1;
        layer_1_weights[375][1] = -1;
        layer_1_weights[376][1] = -2;
        layer_1_weights[377][1] = 0;
        layer_1_weights[378][1] = 1;
        layer_1_weights[379][1] = 0;
        layer_1_weights[380][1] = -1;
        layer_1_weights[381][1] = -2;
        layer_1_weights[382][1] = 0;
        layer_1_weights[383][1] = 0;
        layer_1_weights[384][1] = 1;
        layer_1_weights[385][1] = -1;
        layer_1_weights[386][1] = -2;
        layer_1_weights[387][1] = -1;
        layer_1_weights[388][1] = -2;
        layer_1_weights[389][1] = -1;
        layer_1_weights[390][1] = -1;
        layer_1_weights[391][1] = -1;
        layer_1_weights[392][1] = -1;
        layer_1_weights[393][1] = 1;
        layer_1_weights[394][1] = 4;
        layer_1_weights[395][1] = 0;
        layer_1_weights[396][1] = -1;
        layer_1_weights[397][1] = 0;
        layer_1_weights[398][1] = 0;
        layer_1_weights[399][1] = -3;
        layer_1_weights[400][1] = -3;
        layer_1_weights[401][1] = -1;
        layer_1_weights[402][1] = -1;
        layer_1_weights[403][1] = 0;
        layer_1_weights[404][1] = -1;
        layer_1_weights[405][1] = -1;
        layer_1_weights[406][1] = 1;
        layer_1_weights[407][1] = 2;
        layer_1_weights[408][1] = -1;
        layer_1_weights[409][1] = 1;
        layer_1_weights[410][1] = 1;
        layer_1_weights[411][1] = 1;
        layer_1_weights[412][1] = 0;
        layer_1_weights[413][1] = 1;
        layer_1_weights[414][1] = 0;
        layer_1_weights[415][1] = 0;
        layer_1_weights[416][1] = 0;
        layer_1_weights[417][1] = -7;
        layer_1_weights[418][1] = -3;
        layer_1_weights[419][1] = -2;
        layer_1_weights[420][1] = -2;
        layer_1_weights[421][1] = 1;
        layer_1_weights[422][1] = -3;
        layer_1_weights[423][1] = -2;
        layer_1_weights[424][1] = -3;
        layer_1_weights[425][1] = -2;
        layer_1_weights[426][1] = -2;
        layer_1_weights[427][1] = -3;
        layer_1_weights[428][1] = -2;
        layer_1_weights[429][1] = -2;
        layer_1_weights[430][1] = -1;
        layer_1_weights[431][1] = 0;
        layer_1_weights[432][1] = -1;
        layer_1_weights[433][1] = 1;
        layer_1_weights[434][1] = 0;
        layer_1_weights[435][1] = -1;
        layer_1_weights[436][1] = -1;
        layer_1_weights[437][1] = 0;
        layer_1_weights[438][1] = 2;
        layer_1_weights[439][1] = 1;
        layer_1_weights[440][1] = 0;
        layer_1_weights[441][1] = 1;
        layer_1_weights[442][1] = 0;
        layer_1_weights[443][1] = 0;
        layer_1_weights[444][1] = 0;
        layer_1_weights[445][1] = -3;
        layer_1_weights[446][1] = -2;
        layer_1_weights[447][1] = 0;
        layer_1_weights[448][1] = 2;
        layer_1_weights[449][1] = 3;
        layer_1_weights[450][1] = 0;
        layer_1_weights[451][1] = 1;
        layer_1_weights[452][1] = 0;
        layer_1_weights[453][1] = -1;
        layer_1_weights[454][1] = -2;
        layer_1_weights[455][1] = -2;
        layer_1_weights[456][1] = -2;
        layer_1_weights[457][1] = -2;
        layer_1_weights[458][1] = 0;
        layer_1_weights[459][1] = -1;
        layer_1_weights[460][1] = 1;
        layer_1_weights[461][1] = 0;
        layer_1_weights[462][1] = -1;
        layer_1_weights[463][1] = -1;
        layer_1_weights[464][1] = -1;
        layer_1_weights[465][1] = 1;
        layer_1_weights[466][1] = 2;
        layer_1_weights[467][1] = 2;
        layer_1_weights[468][1] = 0;
        layer_1_weights[469][1] = 0;
        layer_1_weights[470][1] = 0;
        layer_1_weights[471][1] = 0;
        layer_1_weights[472][1] = 1;
        layer_1_weights[473][1] = -6;
        layer_1_weights[474][1] = -4;
        layer_1_weights[475][1] = -1;
        layer_1_weights[476][1] = 1;
        layer_1_weights[477][1] = 2;
        layer_1_weights[478][1] = -2;
        layer_1_weights[479][1] = 4;
        layer_1_weights[480][1] = -1;
        layer_1_weights[481][1] = 0;
        layer_1_weights[482][1] = -2;
        layer_1_weights[483][1] = -1;
        layer_1_weights[484][1] = -1;
        layer_1_weights[485][1] = -2;
        layer_1_weights[486][1] = 0;
        layer_1_weights[487][1] = 0;
        layer_1_weights[488][1] = -1;
        layer_1_weights[489][1] = 0;
        layer_1_weights[490][1] = -2;
        layer_1_weights[491][1] = -1;
        layer_1_weights[492][1] = 1;
        layer_1_weights[493][1] = 1;
        layer_1_weights[494][1] = 1;
        layer_1_weights[495][1] = 2;
        layer_1_weights[496][1] = 0;
        layer_1_weights[497][1] = -2;
        layer_1_weights[498][1] = 1;
        layer_1_weights[499][1] = -2;
        layer_1_weights[500][1] = 1;
        layer_1_weights[501][1] = -1;
        layer_1_weights[502][1] = -1;
        layer_1_weights[503][1] = 1;
        layer_1_weights[504][1] = 3;
        layer_1_weights[505][1] = 1;
        layer_1_weights[506][1] = 1;
        layer_1_weights[507][1] = 1;
        layer_1_weights[508][1] = -2;
        layer_1_weights[509][1] = 1;
        layer_1_weights[510][1] = 0;
        layer_1_weights[511][1] = 0;
        layer_1_weights[512][1] = -2;
        layer_1_weights[513][1] = -1;
        layer_1_weights[514][1] = 0;
        layer_1_weights[515][1] = -1;
        layer_1_weights[516][1] = 0;
        layer_1_weights[517][1] = -1;
        layer_1_weights[518][1] = 0;
        layer_1_weights[519][1] = -1;
        layer_1_weights[520][1] = 1;
        layer_1_weights[521][1] = 1;
        layer_1_weights[522][1] = 1;
        layer_1_weights[523][1] = 1;
        layer_1_weights[524][1] = 1;
        layer_1_weights[525][1] = -1;
        layer_1_weights[526][1] = 1;
        layer_1_weights[527][1] = 0;
        layer_1_weights[528][1] = -1;
        layer_1_weights[529][1] = -1;
        layer_1_weights[530][1] = 3;
        layer_1_weights[531][1] = -4;
        layer_1_weights[532][1] = -1;
        layer_1_weights[533][1] = 2;
        layer_1_weights[534][1] = 2;
        layer_1_weights[535][1] = 1;
        layer_1_weights[536][1] = 0;
        layer_1_weights[537][1] = 0;
        layer_1_weights[538][1] = 1;
        layer_1_weights[539][1] = 0;
        layer_1_weights[540][1] = 0;
        layer_1_weights[541][1] = -1;
        layer_1_weights[542][1] = -1;
        layer_1_weights[543][1] = 0;
        layer_1_weights[544][1] = 1;
        layer_1_weights[545][1] = 0;
        layer_1_weights[546][1] = -1;
        layer_1_weights[547][1] = -1;
        layer_1_weights[548][1] = 1;
        layer_1_weights[549][1] = 0;
        layer_1_weights[550][1] = 0;
        layer_1_weights[551][1] = 0;
        layer_1_weights[552][1] = 0;
        layer_1_weights[553][1] = 0;
        layer_1_weights[554][1] = -1;
        layer_1_weights[555][1] = 0;
        layer_1_weights[556][1] = 0;
        layer_1_weights[557][1] = 0;
        layer_1_weights[558][1] = -3;
        layer_1_weights[559][1] = -3;
        layer_1_weights[560][1] = 0;
        layer_1_weights[561][1] = 2;
        layer_1_weights[562][1] = -3;
        layer_1_weights[563][1] = 0;
        layer_1_weights[564][1] = 0;
        layer_1_weights[565][1] = 0;
        layer_1_weights[566][1] = -1;
        layer_1_weights[567][1] = 1;
        layer_1_weights[568][1] = 1;
        layer_1_weights[569][1] = -1;
        layer_1_weights[570][1] = -1;
        layer_1_weights[571][1] = -1;
        layer_1_weights[572][1] = 0;
        layer_1_weights[573][1] = 0;
        layer_1_weights[574][1] = 1;
        layer_1_weights[575][1] = 0;
        layer_1_weights[576][1] = -1;
        layer_1_weights[577][1] = -1;
        layer_1_weights[578][1] = -1;
        layer_1_weights[579][1] = 1;
        layer_1_weights[580][1] = -1;
        layer_1_weights[581][1] = -1;
        layer_1_weights[582][1] = -1;
        layer_1_weights[583][1] = 1;
        layer_1_weights[584][1] = 1;
        layer_1_weights[585][1] = 1;
        layer_1_weights[586][1] = -4;
        layer_1_weights[587][1] = -2;
        layer_1_weights[588][1] = 0;
        layer_1_weights[589][1] = 1;
        layer_1_weights[590][1] = 1;
        layer_1_weights[591][1] = -2;
        layer_1_weights[592][1] = 0;
        layer_1_weights[593][1] = 1;
        layer_1_weights[594][1] = 1;
        layer_1_weights[595][1] = 0;
        layer_1_weights[596][1] = 1;
        layer_1_weights[597][1] = 1;
        layer_1_weights[598][1] = 0;
        layer_1_weights[599][1] = -1;
        layer_1_weights[600][1] = 1;
        layer_1_weights[601][1] = 1;
        layer_1_weights[602][1] = 1;
        layer_1_weights[603][1] = -1;
        layer_1_weights[604][1] = 0;
        layer_1_weights[605][1] = 0;
        layer_1_weights[606][1] = -1;
        layer_1_weights[607][1] = -2;
        layer_1_weights[608][1] = -1;
        layer_1_weights[609][1] = -1;
        layer_1_weights[610][1] = -2;
        layer_1_weights[611][1] = -2;
        layer_1_weights[612][1] = -2;
        layer_1_weights[613][1] = -2;
        layer_1_weights[614][1] = -3;
        layer_1_weights[615][1] = -1;
        layer_1_weights[616][1] = 0;
        layer_1_weights[617][1] = 2;
        layer_1_weights[618][1] = 0;
        layer_1_weights[619][1] = -1;
        layer_1_weights[620][1] = -1;
        layer_1_weights[621][1] = -1;
        layer_1_weights[622][1] = 2;
        layer_1_weights[623][1] = 2;
        layer_1_weights[624][1] = 1;
        layer_1_weights[625][1] = 1;
        layer_1_weights[626][1] = 0;
        layer_1_weights[627][1] = 1;
        layer_1_weights[628][1] = 1;
        layer_1_weights[629][1] = 1;
        layer_1_weights[630][1] = 2;
        layer_1_weights[631][1] = 0;
        layer_1_weights[632][1] = 0;
        layer_1_weights[633][1] = -1;
        layer_1_weights[634][1] = 0;
        layer_1_weights[635][1] = -3;
        layer_1_weights[636][1] = -2;
        layer_1_weights[637][1] = -4;
        layer_1_weights[638][1] = -2;
        layer_1_weights[639][1] = 1;
        layer_1_weights[640][1] = 0;
        layer_1_weights[641][1] = 1;
        layer_1_weights[642][1] = -1;
        layer_1_weights[643][1] = 0;
        layer_1_weights[644][1] = 0;
        layer_1_weights[645][1] = 0;
        layer_1_weights[646][1] = 1;
        layer_1_weights[647][1] = 1;
        layer_1_weights[648][1] = 2;
        layer_1_weights[649][1] = 1;
        layer_1_weights[650][1] = 1;
        layer_1_weights[651][1] = 2;
        layer_1_weights[652][1] = 0;
        layer_1_weights[653][1] = 0;
        layer_1_weights[654][1] = 0;
        layer_1_weights[655][1] = 0;
        layer_1_weights[656][1] = -1;
        layer_1_weights[657][1] = 0;
        layer_1_weights[658][1] = 0;
        layer_1_weights[659][1] = 1;
        layer_1_weights[660][1] = 1;
        layer_1_weights[661][1] = -1;
        layer_1_weights[662][1] = -1;
        layer_1_weights[663][1] = -3;
        layer_1_weights[664][1] = -1;
        layer_1_weights[665][1] = -1;
        layer_1_weights[666][1] = -2;
        layer_1_weights[667][1] = 2;
        layer_1_weights[668][1] = 3;
        layer_1_weights[669][1] = 2;
        layer_1_weights[670][1] = 0;
        layer_1_weights[671][1] = 0;
        layer_1_weights[672][1] = 0;
        layer_1_weights[673][1] = 0;
        layer_1_weights[674][1] = 1;
        layer_1_weights[675][1] = 3;
        layer_1_weights[676][1] = 4;
        layer_1_weights[677][1] = 5;
        layer_1_weights[678][1] = 1;
        layer_1_weights[679][1] = 1;
        layer_1_weights[680][1] = 0;
        layer_1_weights[681][1] = -2;
        layer_1_weights[682][1] = -1;
        layer_1_weights[683][1] = -1;
        layer_1_weights[684][1] = -1;
        layer_1_weights[685][1] = 1;
        layer_1_weights[686][1] = 1;
        layer_1_weights[687][1] = 1;
        layer_1_weights[688][1] = 0;
        layer_1_weights[689][1] = 1;
        layer_1_weights[690][1] = -1;
        layer_1_weights[691][1] = 0;
        layer_1_weights[692][1] = -1;
        layer_1_weights[693][1] = -1;
        layer_1_weights[694][1] = 0;
        layer_1_weights[695][1] = -1;
        layer_1_weights[696][1] = 2;
        layer_1_weights[697][1] = -5;
        layer_1_weights[698][1] = -2;
        layer_1_weights[699][1] = 0;
        layer_1_weights[700][1] = 0;
        layer_1_weights[701][1] = 0;
        layer_1_weights[702][1] = 3;
        layer_1_weights[703][1] = -1;
        layer_1_weights[704][1] = 1;
        layer_1_weights[705][1] = 2;
        layer_1_weights[706][1] = 2;
        layer_1_weights[707][1] = 1;
        layer_1_weights[708][1] = 3;
        layer_1_weights[709][1] = 1;
        layer_1_weights[710][1] = 3;
        layer_1_weights[711][1] = 4;
        layer_1_weights[712][1] = 5;
        layer_1_weights[713][1] = 2;
        layer_1_weights[714][1] = 3;
        layer_1_weights[715][1] = 2;
        layer_1_weights[716][1] = 4;
        layer_1_weights[717][1] = 4;
        layer_1_weights[718][1] = 2;
        layer_1_weights[719][1] = 4;
        layer_1_weights[720][1] = 4;
        layer_1_weights[721][1] = -1;
        layer_1_weights[722][1] = 2;
        layer_1_weights[723][1] = -1;
        layer_1_weights[724][1] = 2;
        layer_1_weights[725][1] = -1;
        layer_1_weights[726][1] = -2;
        layer_1_weights[727][1] = 0;
        layer_1_weights[728][1] = 0;
        layer_1_weights[729][1] = 1;
        layer_1_weights[730][1] = 0;
        layer_1_weights[731][1] = 2;
        layer_1_weights[732][1] = -2;
        layer_1_weights[733][1] = 0;
        layer_1_weights[734][1] = 1;
        layer_1_weights[735][1] = 5;
        layer_1_weights[736][1] = 6;
        layer_1_weights[737][1] = 4;
        layer_1_weights[738][1] = 5;
        layer_1_weights[739][1] = 6;
        layer_1_weights[740][1] = 7;
        layer_1_weights[741][1] = 6;
        layer_1_weights[742][1] = 7;
        layer_1_weights[743][1] = 7;
        layer_1_weights[744][1] = 5;
        layer_1_weights[745][1] = 7;
        layer_1_weights[746][1] = 5;
        layer_1_weights[747][1] = 5;
        layer_1_weights[748][1] = 6;
        layer_1_weights[749][1] = 9;
        layer_1_weights[750][1] = 5;
        layer_1_weights[751][1] = 0;
        layer_1_weights[752][1] = 0;
        layer_1_weights[753][1] = 2;
        layer_1_weights[754][1] = 0;
        layer_1_weights[755][1] = 0;
        layer_1_weights[756][1] = 0;
        layer_1_weights[757][1] = -1;
        layer_1_weights[758][1] = 0;
        layer_1_weights[759][1] = 1;
        layer_1_weights[760][1] = 1;
        layer_1_weights[761][1] = 3;
        layer_1_weights[762][1] = 2;
        layer_1_weights[763][1] = 4;
        layer_1_weights[764][1] = 4;
        layer_1_weights[765][1] = 5;
        layer_1_weights[766][1] = 5;
        layer_1_weights[767][1] = 5;
        layer_1_weights[768][1] = 5;
        layer_1_weights[769][1] = 7;
        layer_1_weights[770][1] = 7;
        layer_1_weights[771][1] = 5;
        layer_1_weights[772][1] = 3;
        layer_1_weights[773][1] = 7;
        layer_1_weights[774][1] = 4;
        layer_1_weights[775][1] = 3;
        layer_1_weights[776][1] = -1;
        layer_1_weights[777][1] = 3;
        layer_1_weights[778][1] = 3;
        layer_1_weights[779][1] = 3;
        layer_1_weights[780][1] = 1;
        layer_1_weights[781][1] = 0;
        layer_1_weights[782][1] = 1;
        layer_1_weights[783][1] = 1;
        layer_1_weights[0][2] = -1;
        layer_1_weights[1][2] = 0;
        layer_1_weights[2][2] = -1;
        layer_1_weights[3][2] = 1;
        layer_1_weights[4][2] = 0;
        layer_1_weights[5][2] = 0;
        layer_1_weights[6][2] = 1;
        layer_1_weights[7][2] = -1;
        layer_1_weights[8][2] = 1;
        layer_1_weights[9][2] = 0;
        layer_1_weights[10][2] = 0;
        layer_1_weights[11][2] = -1;
        layer_1_weights[12][2] = -1;
        layer_1_weights[13][2] = 0;
        layer_1_weights[14][2] = -1;
        layer_1_weights[15][2] = 0;
        layer_1_weights[16][2] = 1;
        layer_1_weights[17][2] = 0;
        layer_1_weights[18][2] = 0;
        layer_1_weights[19][2] = 0;
        layer_1_weights[20][2] = 0;
        layer_1_weights[21][2] = -1;
        layer_1_weights[22][2] = 1;
        layer_1_weights[23][2] = 1;
        layer_1_weights[24][2] = 0;
        layer_1_weights[25][2] = 0;
        layer_1_weights[26][2] = 0;
        layer_1_weights[27][2] = 0;
        layer_1_weights[28][2] = 0;
        layer_1_weights[29][2] = 0;
        layer_1_weights[30][2] = 0;
        layer_1_weights[31][2] = 0;
        layer_1_weights[32][2] = 0;
        layer_1_weights[33][2] = -1;
        layer_1_weights[34][2] = 1;
        layer_1_weights[35][2] = 0;
        layer_1_weights[36][2] = 0;
        layer_1_weights[37][2] = -2;
        layer_1_weights[38][2] = -1;
        layer_1_weights[39][2] = 0;
        layer_1_weights[40][2] = 0;
        layer_1_weights[41][2] = 2;
        layer_1_weights[42][2] = 3;
        layer_1_weights[43][2] = 3;
        layer_1_weights[44][2] = 1;
        layer_1_weights[45][2] = 1;
        layer_1_weights[46][2] = 1;
        layer_1_weights[47][2] = 0;
        layer_1_weights[48][2] = 0;
        layer_1_weights[49][2] = 0;
        layer_1_weights[50][2] = 0;
        layer_1_weights[51][2] = 0;
        layer_1_weights[52][2] = 0;
        layer_1_weights[53][2] = 0;
        layer_1_weights[54][2] = 0;
        layer_1_weights[55][2] = 1;
        layer_1_weights[56][2] = 0;
        layer_1_weights[57][2] = 0;
        layer_1_weights[58][2] = 0;
        layer_1_weights[59][2] = 0;
        layer_1_weights[60][2] = -1;
        layer_1_weights[61][2] = -1;
        layer_1_weights[62][2] = 1;
        layer_1_weights[63][2] = 1;
        layer_1_weights[64][2] = -1;
        layer_1_weights[65][2] = -1;
        layer_1_weights[66][2] = -1;
        layer_1_weights[67][2] = -1;
        layer_1_weights[68][2] = -1;
        layer_1_weights[69][2] = 2;
        layer_1_weights[70][2] = 5;
        layer_1_weights[71][2] = 4;
        layer_1_weights[72][2] = 5;
        layer_1_weights[73][2] = 5;
        layer_1_weights[74][2] = 5;
        layer_1_weights[75][2] = 4;
        layer_1_weights[76][2] = 4;
        layer_1_weights[77][2] = 2;
        layer_1_weights[78][2] = 3;
        layer_1_weights[79][2] = 2;
        layer_1_weights[80][2] = -1;
        layer_1_weights[81][2] = 0;
        layer_1_weights[82][2] = 0;
        layer_1_weights[83][2] = 0;
        layer_1_weights[84][2] = 0;
        layer_1_weights[85][2] = 0;
        layer_1_weights[86][2] = 0;
        layer_1_weights[87][2] = -3;
        layer_1_weights[88][2] = 0;
        layer_1_weights[89][2] = 0;
        layer_1_weights[90][2] = -4;
        layer_1_weights[91][2] = 1;
        layer_1_weights[92][2] = 0;
        layer_1_weights[93][2] = 2;
        layer_1_weights[94][2] = 0;
        layer_1_weights[95][2] = -2;
        layer_1_weights[96][2] = 1;
        layer_1_weights[97][2] = 3;
        layer_1_weights[98][2] = 2;
        layer_1_weights[99][2] = 4;
        layer_1_weights[100][2] = 0;
        layer_1_weights[101][2] = 0;
        layer_1_weights[102][2] = -1;
        layer_1_weights[103][2] = 3;
        layer_1_weights[104][2] = 2;
        layer_1_weights[105][2] = 2;
        layer_1_weights[106][2] = 0;
        layer_1_weights[107][2] = -3;
        layer_1_weights[108][2] = 5;
        layer_1_weights[109][2] = 3;
        layer_1_weights[110][2] = 3;
        layer_1_weights[111][2] = 0;
        layer_1_weights[112][2] = 1;
        layer_1_weights[113][2] = 1;
        layer_1_weights[114][2] = 0;
        layer_1_weights[115][2] = 1;
        layer_1_weights[116][2] = 0;
        layer_1_weights[117][2] = -1;
        layer_1_weights[118][2] = 0;
        layer_1_weights[119][2] = 0;
        layer_1_weights[120][2] = 0;
        layer_1_weights[121][2] = 0;
        layer_1_weights[122][2] = 1;
        layer_1_weights[123][2] = 0;
        layer_1_weights[124][2] = 0;
        layer_1_weights[125][2] = -1;
        layer_1_weights[126][2] = 0;
        layer_1_weights[127][2] = 0;
        layer_1_weights[128][2] = 0;
        layer_1_weights[129][2] = 1;
        layer_1_weights[130][2] = 1;
        layer_1_weights[131][2] = 1;
        layer_1_weights[132][2] = 1;
        layer_1_weights[133][2] = 2;
        layer_1_weights[134][2] = 2;
        layer_1_weights[135][2] = 3;
        layer_1_weights[136][2] = 1;
        layer_1_weights[137][2] = 6;
        layer_1_weights[138][2] = 3;
        layer_1_weights[139][2] = 0;
        layer_1_weights[140][2] = -1;
        layer_1_weights[141][2] = 0;
        layer_1_weights[142][2] = -2;
        layer_1_weights[143][2] = 1;
        layer_1_weights[144][2] = 2;
        layer_1_weights[145][2] = 4;
        layer_1_weights[146][2] = 0;
        layer_1_weights[147][2] = -1;
        layer_1_weights[148][2] = 1;
        layer_1_weights[149][2] = 0;
        layer_1_weights[150][2] = 0;
        layer_1_weights[151][2] = -1;
        layer_1_weights[152][2] = 1;
        layer_1_weights[153][2] = 2;
        layer_1_weights[154][2] = 2;
        layer_1_weights[155][2] = 0;
        layer_1_weights[156][2] = 0;
        layer_1_weights[157][2] = 1;
        layer_1_weights[158][2] = 2;
        layer_1_weights[159][2] = 2;
        layer_1_weights[160][2] = 1;
        layer_1_weights[161][2] = 2;
        layer_1_weights[162][2] = 1;
        layer_1_weights[163][2] = 3;
        layer_1_weights[164][2] = 3;
        layer_1_weights[165][2] = 2;
        layer_1_weights[166][2] = 5;
        layer_1_weights[167][2] = 3;
        layer_1_weights[168][2] = 1;
        layer_1_weights[169][2] = 0;
        layer_1_weights[170][2] = 0;
        layer_1_weights[171][2] = 2;
        layer_1_weights[172][2] = -2;
        layer_1_weights[173][2] = 3;
        layer_1_weights[174][2] = 1;
        layer_1_weights[175][2] = 1;
        layer_1_weights[176][2] = 0;
        layer_1_weights[177][2] = 2;
        layer_1_weights[178][2] = 1;
        layer_1_weights[179][2] = 0;
        layer_1_weights[180][2] = 1;
        layer_1_weights[181][2] = 1;
        layer_1_weights[182][2] = 1;
        layer_1_weights[183][2] = 1;
        layer_1_weights[184][2] = 1;
        layer_1_weights[185][2] = 2;
        layer_1_weights[186][2] = 1;
        layer_1_weights[187][2] = 1;
        layer_1_weights[188][2] = 2;
        layer_1_weights[189][2] = 1;
        layer_1_weights[190][2] = 2;
        layer_1_weights[191][2] = -2;
        layer_1_weights[192][2] = 0;
        layer_1_weights[193][2] = 3;
        layer_1_weights[194][2] = 1;
        layer_1_weights[195][2] = 2;
        layer_1_weights[196][2] = 0;
        layer_1_weights[197][2] = 3;
        layer_1_weights[198][2] = 3;
        layer_1_weights[199][2] = 1;
        layer_1_weights[200][2] = -1;
        layer_1_weights[201][2] = 1;
        layer_1_weights[202][2] = 2;
        layer_1_weights[203][2] = 1;
        layer_1_weights[204][2] = 1;
        layer_1_weights[205][2] = 2;
        layer_1_weights[206][2] = 2;
        layer_1_weights[207][2] = 1;
        layer_1_weights[208][2] = 2;
        layer_1_weights[209][2] = 2;
        layer_1_weights[210][2] = 1;
        layer_1_weights[211][2] = 3;
        layer_1_weights[212][2] = 2;
        layer_1_weights[213][2] = 2;
        layer_1_weights[214][2] = 1;
        layer_1_weights[215][2] = 1;
        layer_1_weights[216][2] = 2;
        layer_1_weights[217][2] = 1;
        layer_1_weights[218][2] = 1;
        layer_1_weights[219][2] = -2;
        layer_1_weights[220][2] = 1;
        layer_1_weights[221][2] = 0;
        layer_1_weights[222][2] = 3;
        layer_1_weights[223][2] = 0;
        layer_1_weights[224][2] = 0;
        layer_1_weights[225][2] = 1;
        layer_1_weights[226][2] = 2;
        layer_1_weights[227][2] = -2;
        layer_1_weights[228][2] = -2;
        layer_1_weights[229][2] = 1;
        layer_1_weights[230][2] = 1;
        layer_1_weights[231][2] = 0;
        layer_1_weights[232][2] = 2;
        layer_1_weights[233][2] = 2;
        layer_1_weights[234][2] = 2;
        layer_1_weights[235][2] = 2;
        layer_1_weights[236][2] = 4;
        layer_1_weights[237][2] = 2;
        layer_1_weights[238][2] = 3;
        layer_1_weights[239][2] = 2;
        layer_1_weights[240][2] = 0;
        layer_1_weights[241][2] = 0;
        layer_1_weights[242][2] = 0;
        layer_1_weights[243][2] = 0;
        layer_1_weights[244][2] = 0;
        layer_1_weights[245][2] = 0;
        layer_1_weights[246][2] = -2;
        layer_1_weights[247][2] = 0;
        layer_1_weights[248][2] = -1;
        layer_1_weights[249][2] = 0;
        layer_1_weights[250][2] = 5;
        layer_1_weights[251][2] = 1;
        layer_1_weights[252][2] = 1;
        layer_1_weights[253][2] = 2;
        layer_1_weights[254][2] = 4;
        layer_1_weights[255][2] = 0;
        layer_1_weights[256][2] = -1;
        layer_1_weights[257][2] = 1;
        layer_1_weights[258][2] = 0;
        layer_1_weights[259][2] = 1;
        layer_1_weights[260][2] = 2;
        layer_1_weights[261][2] = 2;
        layer_1_weights[262][2] = 2;
        layer_1_weights[263][2] = 1;
        layer_1_weights[264][2] = 3;
        layer_1_weights[265][2] = 3;
        layer_1_weights[266][2] = 2;
        layer_1_weights[267][2] = -1;
        layer_1_weights[268][2] = -2;
        layer_1_weights[269][2] = -3;
        layer_1_weights[270][2] = -2;
        layer_1_weights[271][2] = -2;
        layer_1_weights[272][2] = -2;
        layer_1_weights[273][2] = -2;
        layer_1_weights[274][2] = 0;
        layer_1_weights[275][2] = 1;
        layer_1_weights[276][2] = -3;
        layer_1_weights[277][2] = -1;
        layer_1_weights[278][2] = 2;
        layer_1_weights[279][2] = 2;
        layer_1_weights[280][2] = 1;
        layer_1_weights[281][2] = 4;
        layer_1_weights[282][2] = 4;
        layer_1_weights[283][2] = 1;
        layer_1_weights[284][2] = 1;
        layer_1_weights[285][2] = 0;
        layer_1_weights[286][2] = 1;
        layer_1_weights[287][2] = 0;
        layer_1_weights[288][2] = 2;
        layer_1_weights[289][2] = 0;
        layer_1_weights[290][2] = 1;
        layer_1_weights[291][2] = -1;
        layer_1_weights[292][2] = 1;
        layer_1_weights[293][2] = 0;
        layer_1_weights[294][2] = -1;
        layer_1_weights[295][2] = -3;
        layer_1_weights[296][2] = -4;
        layer_1_weights[297][2] = -3;
        layer_1_weights[298][2] = -3;
        layer_1_weights[299][2] = -3;
        layer_1_weights[300][2] = -3;
        layer_1_weights[301][2] = -2;
        layer_1_weights[302][2] = -2;
        layer_1_weights[303][2] = -4;
        layer_1_weights[304][2] = -3;
        layer_1_weights[305][2] = -4;
        layer_1_weights[306][2] = 5;
        layer_1_weights[307][2] = 2;
        layer_1_weights[308][2] = 2;
        layer_1_weights[309][2] = 4;
        layer_1_weights[310][2] = 3;
        layer_1_weights[311][2] = 0;
        layer_1_weights[312][2] = 1;
        layer_1_weights[313][2] = -1;
        layer_1_weights[314][2] = 0;
        layer_1_weights[315][2] = -1;
        layer_1_weights[316][2] = -1;
        layer_1_weights[317][2] = -1;
        layer_1_weights[318][2] = -1;
        layer_1_weights[319][2] = -1;
        layer_1_weights[320][2] = -2;
        layer_1_weights[321][2] = -2;
        layer_1_weights[322][2] = -3;
        layer_1_weights[323][2] = -4;
        layer_1_weights[324][2] = -1;
        layer_1_weights[325][2] = -2;
        layer_1_weights[326][2] = 0;
        layer_1_weights[327][2] = -1;
        layer_1_weights[328][2] = -2;
        layer_1_weights[329][2] = -3;
        layer_1_weights[330][2] = -2;
        layer_1_weights[331][2] = -2;
        layer_1_weights[332][2] = -5;
        layer_1_weights[333][2] = -6;
        layer_1_weights[334][2] = 3;
        layer_1_weights[335][2] = 2;
        layer_1_weights[336][2] = 1;
        layer_1_weights[337][2] = 1;
        layer_1_weights[338][2] = 1;
        layer_1_weights[339][2] = 1;
        layer_1_weights[340][2] = 2;
        layer_1_weights[341][2] = -1;
        layer_1_weights[342][2] = 0;
        layer_1_weights[343][2] = 0;
        layer_1_weights[344][2] = -1;
        layer_1_weights[345][2] = -1;
        layer_1_weights[346][2] = 0;
        layer_1_weights[347][2] = 0;
        layer_1_weights[348][2] = -1;
        layer_1_weights[349][2] = -4;
        layer_1_weights[350][2] = -3;
        layer_1_weights[351][2] = -1;
        layer_1_weights[352][2] = -1;
        layer_1_weights[353][2] = 0;
        layer_1_weights[354][2] = 1;
        layer_1_weights[355][2] = -1;
        layer_1_weights[356][2] = -1;
        layer_1_weights[357][2] = -1;
        layer_1_weights[358][2] = -2;
        layer_1_weights[359][2] = 0;
        layer_1_weights[360][2] = 0;
        layer_1_weights[361][2] = -8;
        layer_1_weights[362][2] = 0;
        layer_1_weights[363][2] = 1;
        layer_1_weights[364][2] = 0;
        layer_1_weights[365][2] = 0;
        layer_1_weights[366][2] = -1;
        layer_1_weights[367][2] = 1;
        layer_1_weights[368][2] = -2;
        layer_1_weights[369][2] = -1;
        layer_1_weights[370][2] = -2;
        layer_1_weights[371][2] = 0;
        layer_1_weights[372][2] = -2;
        layer_1_weights[373][2] = 0;
        layer_1_weights[374][2] = -1;
        layer_1_weights[375][2] = 0;
        layer_1_weights[376][2] = -2;
        layer_1_weights[377][2] = -1;
        layer_1_weights[378][2] = -1;
        layer_1_weights[379][2] = -2;
        layer_1_weights[380][2] = -1;
        layer_1_weights[381][2] = 0;
        layer_1_weights[382][2] = 1;
        layer_1_weights[383][2] = -1;
        layer_1_weights[384][2] = 1;
        layer_1_weights[385][2] = 1;
        layer_1_weights[386][2] = -1;
        layer_1_weights[387][2] = 1;
        layer_1_weights[388][2] = 0;
        layer_1_weights[389][2] = -5;
        layer_1_weights[390][2] = -1;
        layer_1_weights[391][2] = -1;
        layer_1_weights[392][2] = 3;
        layer_1_weights[393][2] = 1;
        layer_1_weights[394][2] = 3;
        layer_1_weights[395][2] = -2;
        layer_1_weights[396][2] = -2;
        layer_1_weights[397][2] = -1;
        layer_1_weights[398][2] = 1;
        layer_1_weights[399][2] = 0;
        layer_1_weights[400][2] = 1;
        layer_1_weights[401][2] = -1;
        layer_1_weights[402][2] = 0;
        layer_1_weights[403][2] = -1;
        layer_1_weights[404][2] = -2;
        layer_1_weights[405][2] = -1;
        layer_1_weights[406][2] = -1;
        layer_1_weights[407][2] = 0;
        layer_1_weights[408][2] = -1;
        layer_1_weights[409][2] = -1;
        layer_1_weights[410][2] = 0;
        layer_1_weights[411][2] = -2;
        layer_1_weights[412][2] = -1;
        layer_1_weights[413][2] = 1;
        layer_1_weights[414][2] = 0;
        layer_1_weights[415][2] = 3;
        layer_1_weights[416][2] = 2;
        layer_1_weights[417][2] = -5;
        layer_1_weights[418][2] = 0;
        layer_1_weights[419][2] = -1;
        layer_1_weights[420][2] = 3;
        layer_1_weights[421][2] = 0;
        layer_1_weights[422][2] = -2;
        layer_1_weights[423][2] = 0;
        layer_1_weights[424][2] = -2;
        layer_1_weights[425][2] = 0;
        layer_1_weights[426][2] = -2;
        layer_1_weights[427][2] = 0;
        layer_1_weights[428][2] = -2;
        layer_1_weights[429][2] = 0;
        layer_1_weights[430][2] = 0;
        layer_1_weights[431][2] = -1;
        layer_1_weights[432][2] = -1;
        layer_1_weights[433][2] = 0;
        layer_1_weights[434][2] = -1;
        layer_1_weights[435][2] = 0;
        layer_1_weights[436][2] = -2;
        layer_1_weights[437][2] = 0;
        layer_1_weights[438][2] = -2;
        layer_1_weights[439][2] = -2;
        layer_1_weights[440][2] = -1;
        layer_1_weights[441][2] = 1;
        layer_1_weights[442][2] = 1;
        layer_1_weights[443][2] = 1;
        layer_1_weights[444][2] = 3;
        layer_1_weights[445][2] = 3;
        layer_1_weights[446][2] = 3;
        layer_1_weights[447][2] = 1;
        layer_1_weights[448][2] = 1;
        layer_1_weights[449][2] = 0;
        layer_1_weights[450][2] = 2;
        layer_1_weights[451][2] = -1;
        layer_1_weights[452][2] = -1;
        layer_1_weights[453][2] = 0;
        layer_1_weights[454][2] = -1;
        layer_1_weights[455][2] = -1;
        layer_1_weights[456][2] = 0;
        layer_1_weights[457][2] = 0;
        layer_1_weights[458][2] = 0;
        layer_1_weights[459][2] = 1;
        layer_1_weights[460][2] = -1;
        layer_1_weights[461][2] = -1;
        layer_1_weights[462][2] = -1;
        layer_1_weights[463][2] = 0;
        layer_1_weights[464][2] = -2;
        layer_1_weights[465][2] = -1;
        layer_1_weights[466][2] = 0;
        layer_1_weights[467][2] = -1;
        layer_1_weights[468][2] = 0;
        layer_1_weights[469][2] = 1;
        layer_1_weights[470][2] = 1;
        layer_1_weights[471][2] = 2;
        layer_1_weights[472][2] = -1;
        layer_1_weights[473][2] = 1;
        layer_1_weights[474][2] = -2;
        layer_1_weights[475][2] = 1;
        layer_1_weights[476][2] = -1;
        layer_1_weights[477][2] = 0;
        layer_1_weights[478][2] = -1;
        layer_1_weights[479][2] = 4;
        layer_1_weights[480][2] = 1;
        layer_1_weights[481][2] = -3;
        layer_1_weights[482][2] = -2;
        layer_1_weights[483][2] = -1;
        layer_1_weights[484][2] = -2;
        layer_1_weights[485][2] = -2;
        layer_1_weights[486][2] = -1;
        layer_1_weights[487][2] = -1;
        layer_1_weights[488][2] = -1;
        layer_1_weights[489][2] = -2;
        layer_1_weights[490][2] = -2;
        layer_1_weights[491][2] = -2;
        layer_1_weights[492][2] = -2;
        layer_1_weights[493][2] = -2;
        layer_1_weights[494][2] = -1;
        layer_1_weights[495][2] = 1;
        layer_1_weights[496][2] = 1;
        layer_1_weights[497][2] = 1;
        layer_1_weights[498][2] = 0;
        layer_1_weights[499][2] = 2;
        layer_1_weights[500][2] = 1;
        layer_1_weights[501][2] = 1;
        layer_1_weights[502][2] = -3;
        layer_1_weights[503][2] = -3;
        layer_1_weights[504][2] = 1;
        layer_1_weights[505][2] = -1;
        layer_1_weights[506][2] = -1;
        layer_1_weights[507][2] = 3;
        layer_1_weights[508][2] = 1;
        layer_1_weights[509][2] = -3;
        layer_1_weights[510][2] = -1;
        layer_1_weights[511][2] = -1;
        layer_1_weights[512][2] = -1;
        layer_1_weights[513][2] = -2;
        layer_1_weights[514][2] = -2;
        layer_1_weights[515][2] = -2;
        layer_1_weights[516][2] = -4;
        layer_1_weights[517][2] = -4;
        layer_1_weights[518][2] = -2;
        layer_1_weights[519][2] = -1;
        layer_1_weights[520][2] = 0;
        layer_1_weights[521][2] = 0;
        layer_1_weights[522][2] = -1;
        layer_1_weights[523][2] = 0;
        layer_1_weights[524][2] = 0;
        layer_1_weights[525][2] = 2;
        layer_1_weights[526][2] = 1;
        layer_1_weights[527][2] = 1;
        layer_1_weights[528][2] = -2;
        layer_1_weights[529][2] = 1;
        layer_1_weights[530][2] = -3;
        layer_1_weights[531][2] = -2;
        layer_1_weights[532][2] = -1;
        layer_1_weights[533][2] = 0;
        layer_1_weights[534][2] = 4;
        layer_1_weights[535][2] = 2;
        layer_1_weights[536][2] = 1;
        layer_1_weights[537][2] = -2;
        layer_1_weights[538][2] = 0;
        layer_1_weights[539][2] = -2;
        layer_1_weights[540][2] = -1;
        layer_1_weights[541][2] = -2;
        layer_1_weights[542][2] = -3;
        layer_1_weights[543][2] = -2;
        layer_1_weights[544][2] = -1;
        layer_1_weights[545][2] = -3;
        layer_1_weights[546][2] = 0;
        layer_1_weights[547][2] = 1;
        layer_1_weights[548][2] = 0;
        layer_1_weights[549][2] = 0;
        layer_1_weights[550][2] = 0;
        layer_1_weights[551][2] = 1;
        layer_1_weights[552][2] = 1;
        layer_1_weights[553][2] = 1;
        layer_1_weights[554][2] = 0;
        layer_1_weights[555][2] = 0;
        layer_1_weights[556][2] = 0;
        layer_1_weights[557][2] = 2;
        layer_1_weights[558][2] = -4;
        layer_1_weights[559][2] = -2;
        layer_1_weights[560][2] = 0;
        layer_1_weights[561][2] = 1;
        layer_1_weights[562][2] = 1;
        layer_1_weights[563][2] = 2;
        layer_1_weights[564][2] = 0;
        layer_1_weights[565][2] = 0;
        layer_1_weights[566][2] = 0;
        layer_1_weights[567][2] = 0;
        layer_1_weights[568][2] = -1;
        layer_1_weights[569][2] = -1;
        layer_1_weights[570][2] = -1;
        layer_1_weights[571][2] = 0;
        layer_1_weights[572][2] = 0;
        layer_1_weights[573][2] = 1;
        layer_1_weights[574][2] = 2;
        layer_1_weights[575][2] = 1;
        layer_1_weights[576][2] = 2;
        layer_1_weights[577][2] = 0;
        layer_1_weights[578][2] = 0;
        layer_1_weights[579][2] = 0;
        layer_1_weights[580][2] = 1;
        layer_1_weights[581][2] = 0;
        layer_1_weights[582][2] = 1;
        layer_1_weights[583][2] = -1;
        layer_1_weights[584][2] = -1;
        layer_1_weights[585][2] = 0;
        layer_1_weights[586][2] = 0;
        layer_1_weights[587][2] = 1;
        layer_1_weights[588][2] = 0;
        layer_1_weights[589][2] = 0;
        layer_1_weights[590][2] = -2;
        layer_1_weights[591][2] = 3;
        layer_1_weights[592][2] = 2;
        layer_1_weights[593][2] = 0;
        layer_1_weights[594][2] = 0;
        layer_1_weights[595][2] = 0;
        layer_1_weights[596][2] = 1;
        layer_1_weights[597][2] = 1;
        layer_1_weights[598][2] = 1;
        layer_1_weights[599][2] = 2;
        layer_1_weights[600][2] = 2;
        layer_1_weights[601][2] = 2;
        layer_1_weights[602][2] = 3;
        layer_1_weights[603][2] = 3;
        layer_1_weights[604][2] = 2;
        layer_1_weights[605][2] = 0;
        layer_1_weights[606][2] = 1;
        layer_1_weights[607][2] = 0;
        layer_1_weights[608][2] = 2;
        layer_1_weights[609][2] = 1;
        layer_1_weights[610][2] = 2;
        layer_1_weights[611][2] = 0;
        layer_1_weights[612][2] = -1;
        layer_1_weights[613][2] = 0;
        layer_1_weights[614][2] = 1;
        layer_1_weights[615][2] = 1;
        layer_1_weights[616][2] = -1;
        layer_1_weights[617][2] = -1;
        layer_1_weights[618][2] = -2;
        layer_1_weights[619][2] = 1;
        layer_1_weights[620][2] = 0;
        layer_1_weights[621][2] = 2;
        layer_1_weights[622][2] = 0;
        layer_1_weights[623][2] = 1;
        layer_1_weights[624][2] = 2;
        layer_1_weights[625][2] = 1;
        layer_1_weights[626][2] = 0;
        layer_1_weights[627][2] = 2;
        layer_1_weights[628][2] = 2;
        layer_1_weights[629][2] = 2;
        layer_1_weights[630][2] = 2;
        layer_1_weights[631][2] = 1;
        layer_1_weights[632][2] = 2;
        layer_1_weights[633][2] = 1;
        layer_1_weights[634][2] = 2;
        layer_1_weights[635][2] = 0;
        layer_1_weights[636][2] = 3;
        layer_1_weights[637][2] = 0;
        layer_1_weights[638][2] = 1;
        layer_1_weights[639][2] = 2;
        layer_1_weights[640][2] = 0;
        layer_1_weights[641][2] = 1;
        layer_1_weights[642][2] = -2;
        layer_1_weights[643][2] = 2;
        layer_1_weights[644][2] = 0;
        layer_1_weights[645][2] = 0;
        layer_1_weights[646][2] = 2;
        layer_1_weights[647][2] = 2;
        layer_1_weights[648][2] = 4;
        layer_1_weights[649][2] = 1;
        layer_1_weights[650][2] = 1;
        layer_1_weights[651][2] = -1;
        layer_1_weights[652][2] = 2;
        layer_1_weights[653][2] = 1;
        layer_1_weights[654][2] = 1;
        layer_1_weights[655][2] = 1;
        layer_1_weights[656][2] = 0;
        layer_1_weights[657][2] = 1;
        layer_1_weights[658][2] = -1;
        layer_1_weights[659][2] = 1;
        layer_1_weights[660][2] = 1;
        layer_1_weights[661][2] = 1;
        layer_1_weights[662][2] = 2;
        layer_1_weights[663][2] = 2;
        layer_1_weights[664][2] = 0;
        layer_1_weights[665][2] = 1;
        layer_1_weights[666][2] = -2;
        layer_1_weights[667][2] = 0;
        layer_1_weights[668][2] = -3;
        layer_1_weights[669][2] = -2;
        layer_1_weights[670][2] = 0;
        layer_1_weights[671][2] = -1;
        layer_1_weights[672][2] = 0;
        layer_1_weights[673][2] = 0;
        layer_1_weights[674][2] = -2;
        layer_1_weights[675][2] = 4;
        layer_1_weights[676][2] = 5;
        layer_1_weights[677][2] = 3;
        layer_1_weights[678][2] = 2;
        layer_1_weights[679][2] = 3;
        layer_1_weights[680][2] = 1;
        layer_1_weights[681][2] = 2;
        layer_1_weights[682][2] = 2;
        layer_1_weights[683][2] = 2;
        layer_1_weights[684][2] = 1;
        layer_1_weights[685][2] = 1;
        layer_1_weights[686][2] = 2;
        layer_1_weights[687][2] = 1;
        layer_1_weights[688][2] = 1;
        layer_1_weights[689][2] = 1;
        layer_1_weights[690][2] = 2;
        layer_1_weights[691][2] = 1;
        layer_1_weights[692][2] = 1;
        layer_1_weights[693][2] = -1;
        layer_1_weights[694][2] = 0;
        layer_1_weights[695][2] = -1;
        layer_1_weights[696][2] = 1;
        layer_1_weights[697][2] = -3;
        layer_1_weights[698][2] = 0;
        layer_1_weights[699][2] = -1;
        layer_1_weights[700][2] = 0;
        layer_1_weights[701][2] = 0;
        layer_1_weights[702][2] = -2;
        layer_1_weights[703][2] = 3;
        layer_1_weights[704][2] = 5;
        layer_1_weights[705][2] = 2;
        layer_1_weights[706][2] = 2;
        layer_1_weights[707][2] = 7;
        layer_1_weights[708][2] = 5;
        layer_1_weights[709][2] = 6;
        layer_1_weights[710][2] = 4;
        layer_1_weights[711][2] = 3;
        layer_1_weights[712][2] = 2;
        layer_1_weights[713][2] = 2;
        layer_1_weights[714][2] = -1;
        layer_1_weights[715][2] = 0;
        layer_1_weights[716][2] = 1;
        layer_1_weights[717][2] = 2;
        layer_1_weights[718][2] = 1;
        layer_1_weights[719][2] = -1;
        layer_1_weights[720][2] = 1;
        layer_1_weights[721][2] = 1;
        layer_1_weights[722][2] = 3;
        layer_1_weights[723][2] = 0;
        layer_1_weights[724][2] = 2;
        layer_1_weights[725][2] = -2;
        layer_1_weights[726][2] = 0;
        layer_1_weights[727][2] = -1;
        layer_1_weights[728][2] = 1;
        layer_1_weights[729][2] = -1;
        layer_1_weights[730][2] = 0;
        layer_1_weights[731][2] = -1;
        layer_1_weights[732][2] = 2;
        layer_1_weights[733][2] = 1;
        layer_1_weights[734][2] = 3;
        layer_1_weights[735][2] = 3;
        layer_1_weights[736][2] = 3;
        layer_1_weights[737][2] = 2;
        layer_1_weights[738][2] = 2;
        layer_1_weights[739][2] = 2;
        layer_1_weights[740][2] = 0;
        layer_1_weights[741][2] = 4;
        layer_1_weights[742][2] = 2;
        layer_1_weights[743][2] = 4;
        layer_1_weights[744][2] = 1;
        layer_1_weights[745][2] = 1;
        layer_1_weights[746][2] = 1;
        layer_1_weights[747][2] = 3;
        layer_1_weights[748][2] = 1;
        layer_1_weights[749][2] = 1;
        layer_1_weights[750][2] = 4;
        layer_1_weights[751][2] = -1;
        layer_1_weights[752][2] = 0;
        layer_1_weights[753][2] = 1;
        layer_1_weights[754][2] = 1;
        layer_1_weights[755][2] = -1;
        layer_1_weights[756][2] = -1;
        layer_1_weights[757][2] = 0;
        layer_1_weights[758][2] = 0;
        layer_1_weights[759][2] = 0;
        layer_1_weights[760][2] = 0;
        layer_1_weights[761][2] = 3;
        layer_1_weights[762][2] = 4;
        layer_1_weights[763][2] = 6;
        layer_1_weights[764][2] = 6;
        layer_1_weights[765][2] = 3;
        layer_1_weights[766][2] = 5;
        layer_1_weights[767][2] = 6;
        layer_1_weights[768][2] = 7;
        layer_1_weights[769][2] = 5;
        layer_1_weights[770][2] = 5;
        layer_1_weights[771][2] = 0;
        layer_1_weights[772][2] = 0;
        layer_1_weights[773][2] = 6;
        layer_1_weights[774][2] = 0;
        layer_1_weights[775][2] = -1;
        layer_1_weights[776][2] = 0;
        layer_1_weights[777][2] = 1;
        layer_1_weights[778][2] = 0;
        layer_1_weights[779][2] = 0;
        layer_1_weights[780][2] = 1;
        layer_1_weights[781][2] = 0;
        layer_1_weights[782][2] = 0;
        layer_1_weights[783][2] = 0;
        layer_1_weights[0][3] = -1;
        layer_1_weights[1][3] = -1;
        layer_1_weights[2][3] = 0;
        layer_1_weights[3][3] = 0;
        layer_1_weights[4][3] = 0;
        layer_1_weights[5][3] = 0;
        layer_1_weights[6][3] = 0;
        layer_1_weights[7][3] = 1;
        layer_1_weights[8][3] = 1;
        layer_1_weights[9][3] = 0;
        layer_1_weights[10][3] = 0;
        layer_1_weights[11][3] = 1;
        layer_1_weights[12][3] = -2;
        layer_1_weights[13][3] = 0;
        layer_1_weights[14][3] = 2;
        layer_1_weights[15][3] = 0;
        layer_1_weights[16][3] = 0;
        layer_1_weights[17][3] = -1;
        layer_1_weights[18][3] = 0;
        layer_1_weights[19][3] = 1;
        layer_1_weights[20][3] = 0;
        layer_1_weights[21][3] = 0;
        layer_1_weights[22][3] = 0;
        layer_1_weights[23][3] = 1;
        layer_1_weights[24][3] = 0;
        layer_1_weights[25][3] = 0;
        layer_1_weights[26][3] = 0;
        layer_1_weights[27][3] = 0;
        layer_1_weights[28][3] = 0;
        layer_1_weights[29][3] = 0;
        layer_1_weights[30][3] = -1;
        layer_1_weights[31][3] = 0;
        layer_1_weights[32][3] = -1;
        layer_1_weights[33][3] = -2;
        layer_1_weights[34][3] = -3;
        layer_1_weights[35][3] = -3;
        layer_1_weights[36][3] = -3;
        layer_1_weights[37][3] = -4;
        layer_1_weights[38][3] = -6;
        layer_1_weights[39][3] = 0;
        layer_1_weights[40][3] = -3;
        layer_1_weights[41][3] = -3;
        layer_1_weights[42][3] = 1;
        layer_1_weights[43][3] = -4;
        layer_1_weights[44][3] = -2;
        layer_1_weights[45][3] = -4;
        layer_1_weights[46][3] = -5;
        layer_1_weights[47][3] = -5;
        layer_1_weights[48][3] = -3;
        layer_1_weights[49][3] = -3;
        layer_1_weights[50][3] = -2;
        layer_1_weights[51][3] = -2;
        layer_1_weights[52][3] = 1;
        layer_1_weights[53][3] = 0;
        layer_1_weights[54][3] = 0;
        layer_1_weights[55][3] = 0;
        layer_1_weights[56][3] = 0;
        layer_1_weights[57][3] = 0;
        layer_1_weights[58][3] = -1;
        layer_1_weights[59][3] = 0;
        layer_1_weights[60][3] = -2;
        layer_1_weights[61][3] = -1;
        layer_1_weights[62][3] = -3;
        layer_1_weights[63][3] = -7;
        layer_1_weights[64][3] = -3;
        layer_1_weights[65][3] = -3;
        layer_1_weights[66][3] = -6;
        layer_1_weights[67][3] = -8;
        layer_1_weights[68][3] = -5;
        layer_1_weights[69][3] = -1;
        layer_1_weights[70][3] = 0;
        layer_1_weights[71][3] = -2;
        layer_1_weights[72][3] = -2;
        layer_1_weights[73][3] = -1;
        layer_1_weights[74][3] = -4;
        layer_1_weights[75][3] = -1;
        layer_1_weights[76][3] = -5;
        layer_1_weights[77][3] = -4;
        layer_1_weights[78][3] = -3;
        layer_1_weights[79][3] = -5;
        layer_1_weights[80][3] = -3;
        layer_1_weights[81][3] = -1;
        layer_1_weights[82][3] = 0;
        layer_1_weights[83][3] = 0;
        layer_1_weights[84][3] = 0;
        layer_1_weights[85][3] = 0;
        layer_1_weights[86][3] = -1;
        layer_1_weights[87][3] = -3;
        layer_1_weights[88][3] = 1;
        layer_1_weights[89][3] = -4;
        layer_1_weights[90][3] = -3;
        layer_1_weights[91][3] = -5;
        layer_1_weights[92][3] = -3;
        layer_1_weights[93][3] = -1;
        layer_1_weights[94][3] = 0;
        layer_1_weights[95][3] = 0;
        layer_1_weights[96][3] = -2;
        layer_1_weights[97][3] = -3;
        layer_1_weights[98][3] = 0;
        layer_1_weights[99][3] = -2;
        layer_1_weights[100][3] = -3;
        layer_1_weights[101][3] = -2;
        layer_1_weights[102][3] = -2;
        layer_1_weights[103][3] = -1;
        layer_1_weights[104][3] = 1;
        layer_1_weights[105][3] = 2;
        layer_1_weights[106][3] = 0;
        layer_1_weights[107][3] = -3;
        layer_1_weights[108][3] = -4;
        layer_1_weights[109][3] = -2;
        layer_1_weights[110][3] = 0;
        layer_1_weights[111][3] = 0;
        layer_1_weights[112][3] = 1;
        layer_1_weights[113][3] = -2;
        layer_1_weights[114][3] = 0;
        layer_1_weights[115][3] = -2;
        layer_1_weights[116][3] = -3;
        layer_1_weights[117][3] = -5;
        layer_1_weights[118][3] = -1;
        layer_1_weights[119][3] = 1;
        layer_1_weights[120][3] = 0;
        layer_1_weights[121][3] = 1;
        layer_1_weights[122][3] = -2;
        layer_1_weights[123][3] = 1;
        layer_1_weights[124][3] = 0;
        layer_1_weights[125][3] = 2;
        layer_1_weights[126][3] = 0;
        layer_1_weights[127][3] = 1;
        layer_1_weights[128][3] = 0;
        layer_1_weights[129][3] = 1;
        layer_1_weights[130][3] = 2;
        layer_1_weights[131][3] = 0;
        layer_1_weights[132][3] = -2;
        layer_1_weights[133][3] = -5;
        layer_1_weights[134][3] = -2;
        layer_1_weights[135][3] = -1;
        layer_1_weights[136][3] = 0;
        layer_1_weights[137][3] = 1;
        layer_1_weights[138][3] = -2;
        layer_1_weights[139][3] = -3;
        layer_1_weights[140][3] = 0;
        layer_1_weights[141][3] = 1;
        layer_1_weights[142][3] = -2;
        layer_1_weights[143][3] = 2;
        layer_1_weights[144][3] = -4;
        layer_1_weights[145][3] = 0;
        layer_1_weights[146][3] = 1;
        layer_1_weights[147][3] = 1;
        layer_1_weights[148][3] = 3;
        layer_1_weights[149][3] = 2;
        layer_1_weights[150][3] = 2;
        layer_1_weights[151][3] = -2;
        layer_1_weights[152][3] = -1;
        layer_1_weights[153][3] = 0;
        layer_1_weights[154][3] = -1;
        layer_1_weights[155][3] = -1;
        layer_1_weights[156][3] = 0;
        layer_1_weights[157][3] = -2;
        layer_1_weights[158][3] = -2;
        layer_1_weights[159][3] = -3;
        layer_1_weights[160][3] = -3;
        layer_1_weights[161][3] = -2;
        layer_1_weights[162][3] = -1;
        layer_1_weights[163][3] = -2;
        layer_1_weights[164][3] = -2;
        layer_1_weights[165][3] = 1;
        layer_1_weights[166][3] = -1;
        layer_1_weights[167][3] = -1;
        layer_1_weights[168][3] = 0;
        layer_1_weights[169][3] = 1;
        layer_1_weights[170][3] = 1;
        layer_1_weights[171][3] = -1;
        layer_1_weights[172][3] = 1;
        layer_1_weights[173][3] = 2;
        layer_1_weights[174][3] = 1;
        layer_1_weights[175][3] = 2;
        layer_1_weights[176][3] = 1;
        layer_1_weights[177][3] = 1;
        layer_1_weights[178][3] = 0;
        layer_1_weights[179][3] = 1;
        layer_1_weights[180][3] = 0;
        layer_1_weights[181][3] = -1;
        layer_1_weights[182][3] = 0;
        layer_1_weights[183][3] = -3;
        layer_1_weights[184][3] = -2;
        layer_1_weights[185][3] = -1;
        layer_1_weights[186][3] = -3;
        layer_1_weights[187][3] = -1;
        layer_1_weights[188][3] = -2;
        layer_1_weights[189][3] = -1;
        layer_1_weights[190][3] = 0;
        layer_1_weights[191][3] = 1;
        layer_1_weights[192][3] = 0;
        layer_1_weights[193][3] = 1;
        layer_1_weights[194][3] = 2;
        layer_1_weights[195][3] = -1;
        layer_1_weights[196][3] = 1;
        layer_1_weights[197][3] = -2;
        layer_1_weights[198][3] = 0;
        layer_1_weights[199][3] = 2;
        layer_1_weights[200][3] = -1;
        layer_1_weights[201][3] = 2;
        layer_1_weights[202][3] = 3;
        layer_1_weights[203][3] = 1;
        layer_1_weights[204][3] = 2;
        layer_1_weights[205][3] = 1;
        layer_1_weights[206][3] = 1;
        layer_1_weights[207][3] = 0;
        layer_1_weights[208][3] = -1;
        layer_1_weights[209][3] = -2;
        layer_1_weights[210][3] = -1;
        layer_1_weights[211][3] = -2;
        layer_1_weights[212][3] = -1;
        layer_1_weights[213][3] = 0;
        layer_1_weights[214][3] = 0;
        layer_1_weights[215][3] = 0;
        layer_1_weights[216][3] = 2;
        layer_1_weights[217][3] = 2;
        layer_1_weights[218][3] = 3;
        layer_1_weights[219][3] = 3;
        layer_1_weights[220][3] = 3;
        layer_1_weights[221][3] = 3;
        layer_1_weights[222][3] = 5;
        layer_1_weights[223][3] = -1;
        layer_1_weights[224][3] = 0;
        layer_1_weights[225][3] = 2;
        layer_1_weights[226][3] = 4;
        layer_1_weights[227][3] = 3;
        layer_1_weights[228][3] = -1;
        layer_1_weights[229][3] = 1;
        layer_1_weights[230][3] = 0;
        layer_1_weights[231][3] = 1;
        layer_1_weights[232][3] = 1;
        layer_1_weights[233][3] = 1;
        layer_1_weights[234][3] = 0;
        layer_1_weights[235][3] = -1;
        layer_1_weights[236][3] = 0;
        layer_1_weights[237][3] = -1;
        layer_1_weights[238][3] = 0;
        layer_1_weights[239][3] = 0;
        layer_1_weights[240][3] = -1;
        layer_1_weights[241][3] = 1;
        layer_1_weights[242][3] = 0;
        layer_1_weights[243][3] = 0;
        layer_1_weights[244][3] = 1;
        layer_1_weights[245][3] = 2;
        layer_1_weights[246][3] = 0;
        layer_1_weights[247][3] = 1;
        layer_1_weights[248][3] = 4;
        layer_1_weights[249][3] = 5;
        layer_1_weights[250][3] = 0;
        layer_1_weights[251][3] = 2;
        layer_1_weights[252][3] = 2;
        layer_1_weights[253][3] = 3;
        layer_1_weights[254][3] = 0;
        layer_1_weights[255][3] = 1;
        layer_1_weights[256][3] = -1;
        layer_1_weights[257][3] = 2;
        layer_1_weights[258][3] = -1;
        layer_1_weights[259][3] = 0;
        layer_1_weights[260][3] = 1;
        layer_1_weights[261][3] = 0;
        layer_1_weights[262][3] = 1;
        layer_1_weights[263][3] = 2;
        layer_1_weights[264][3] = -1;
        layer_1_weights[265][3] = -2;
        layer_1_weights[266][3] = -1;
        layer_1_weights[267][3] = 0;
        layer_1_weights[268][3] = 0;
        layer_1_weights[269][3] = 2;
        layer_1_weights[270][3] = 2;
        layer_1_weights[271][3] = 2;
        layer_1_weights[272][3] = 1;
        layer_1_weights[273][3] = 1;
        layer_1_weights[274][3] = 1;
        layer_1_weights[275][3] = 2;
        layer_1_weights[276][3] = 5;
        layer_1_weights[277][3] = 6;
        layer_1_weights[278][3] = 3;
        layer_1_weights[279][3] = 0;
        layer_1_weights[280][3] = 2;
        layer_1_weights[281][3] = 3;
        layer_1_weights[282][3] = 1;
        layer_1_weights[283][3] = -2;
        layer_1_weights[284][3] = 2;
        layer_1_weights[285][3] = 1;
        layer_1_weights[286][3] = 1;
        layer_1_weights[287][3] = 1;
        layer_1_weights[288][3] = 0;
        layer_1_weights[289][3] = 2;
        layer_1_weights[290][3] = 1;
        layer_1_weights[291][3] = 1;
        layer_1_weights[292][3] = 0;
        layer_1_weights[293][3] = -2;
        layer_1_weights[294][3] = -2;
        layer_1_weights[295][3] = 1;
        layer_1_weights[296][3] = 0;
        layer_1_weights[297][3] = 1;
        layer_1_weights[298][3] = 1;
        layer_1_weights[299][3] = 2;
        layer_1_weights[300][3] = 0;
        layer_1_weights[301][3] = 1;
        layer_1_weights[302][3] = -1;
        layer_1_weights[303][3] = -1;
        layer_1_weights[304][3] = 2;
        layer_1_weights[305][3] = 3;
        layer_1_weights[306][3] = 5;
        layer_1_weights[307][3] = -1;
        layer_1_weights[308][3] = 4;
        layer_1_weights[309][3] = 2;
        layer_1_weights[310][3] = -1;
        layer_1_weights[311][3] = 1;
        layer_1_weights[312][3] = 0;
        layer_1_weights[313][3] = -1;
        layer_1_weights[314][3] = 1;
        layer_1_weights[315][3] = 0;
        layer_1_weights[316][3] = 1;
        layer_1_weights[317][3] = 1;
        layer_1_weights[318][3] = 2;
        layer_1_weights[319][3] = 2;
        layer_1_weights[320][3] = 0;
        layer_1_weights[321][3] = -1;
        layer_1_weights[322][3] = -2;
        layer_1_weights[323][3] = -1;
        layer_1_weights[324][3] = 0;
        layer_1_weights[325][3] = -1;
        layer_1_weights[326][3] = 1;
        layer_1_weights[327][3] = 0;
        layer_1_weights[328][3] = -2;
        layer_1_weights[329][3] = -1;
        layer_1_weights[330][3] = -3;
        layer_1_weights[331][3] = -2;
        layer_1_weights[332][3] = 0;
        layer_1_weights[333][3] = 2;
        layer_1_weights[334][3] = 1;
        layer_1_weights[335][3] = 1;
        layer_1_weights[336][3] = 2;
        layer_1_weights[337][3] = 6;
        layer_1_weights[338][3] = 3;
        layer_1_weights[339][3] = -1;
        layer_1_weights[340][3] = -2;
        layer_1_weights[341][3] = 0;
        layer_1_weights[342][3] = 1;
        layer_1_weights[343][3] = 1;
        layer_1_weights[344][3] = 1;
        layer_1_weights[345][3] = 1;
        layer_1_weights[346][3] = 2;
        layer_1_weights[347][3] = 3;
        layer_1_weights[348][3] = 1;
        layer_1_weights[349][3] = -1;
        layer_1_weights[350][3] = -3;
        layer_1_weights[351][3] = -2;
        layer_1_weights[352][3] = 1;
        layer_1_weights[353][3] = 0;
        layer_1_weights[354][3] = -1;
        layer_1_weights[355][3] = 0;
        layer_1_weights[356][3] = -1;
        layer_1_weights[357][3] = -1;
        layer_1_weights[358][3] = -1;
        layer_1_weights[359][3] = -4;
        layer_1_weights[360][3] = -4;
        layer_1_weights[361][3] = 0;
        layer_1_weights[362][3] = 4;
        layer_1_weights[363][3] = -2;
        layer_1_weights[364][3] = 0;
        layer_1_weights[365][3] = 4;
        layer_1_weights[366][3] = 4;
        layer_1_weights[367][3] = 1;
        layer_1_weights[368][3] = -1;
        layer_1_weights[369][3] = 2;
        layer_1_weights[370][3] = 0;
        layer_1_weights[371][3] = 1;
        layer_1_weights[372][3] = 1;
        layer_1_weights[373][3] = 2;
        layer_1_weights[374][3] = 3;
        layer_1_weights[375][3] = 2;
        layer_1_weights[376][3] = 1;
        layer_1_weights[377][3] = -3;
        layer_1_weights[378][3] = -2;
        layer_1_weights[379][3] = 0;
        layer_1_weights[380][3] = -1;
        layer_1_weights[381][3] = -2;
        layer_1_weights[382][3] = 1;
        layer_1_weights[383][3] = -2;
        layer_1_weights[384][3] = 0;
        layer_1_weights[385][3] = 0;
        layer_1_weights[386][3] = 1;
        layer_1_weights[387][3] = -4;
        layer_1_weights[388][3] = -2;
        layer_1_weights[389][3] = 2;
        layer_1_weights[390][3] = 2;
        layer_1_weights[391][3] = -4;
        layer_1_weights[392][3] = 2;
        layer_1_weights[393][3] = -1;
        layer_1_weights[394][3] = 5;
        layer_1_weights[395][3] = 2;
        layer_1_weights[396][3] = -1;
        layer_1_weights[397][3] = 1;
        layer_1_weights[398][3] = 2;
        layer_1_weights[399][3] = 2;
        layer_1_weights[400][3] = 1;
        layer_1_weights[401][3] = 1;
        layer_1_weights[402][3] = 2;
        layer_1_weights[403][3] = 3;
        layer_1_weights[404][3] = 0;
        layer_1_weights[405][3] = -2;
        layer_1_weights[406][3] = -1;
        layer_1_weights[407][3] = -1;
        layer_1_weights[408][3] = 0;
        layer_1_weights[409][3] = 0;
        layer_1_weights[410][3] = 1;
        layer_1_weights[411][3] = 1;
        layer_1_weights[412][3] = 0;
        layer_1_weights[413][3] = 0;
        layer_1_weights[414][3] = 1;
        layer_1_weights[415][3] = 2;
        layer_1_weights[416][3] = 3;
        layer_1_weights[417][3] = 0;
        layer_1_weights[418][3] = -1;
        layer_1_weights[419][3] = 0;
        layer_1_weights[420][3] = 1;
        layer_1_weights[421][3] = -1;
        layer_1_weights[422][3] = 2;
        layer_1_weights[423][3] = 1;
        layer_1_weights[424][3] = 0;
        layer_1_weights[425][3] = 1;
        layer_1_weights[426][3] = 0;
        layer_1_weights[427][3] = 2;
        layer_1_weights[428][3] = 0;
        layer_1_weights[429][3] = 0;
        layer_1_weights[430][3] = 0;
        layer_1_weights[431][3] = 1;
        layer_1_weights[432][3] = -2;
        layer_1_weights[433][3] = -3;
        layer_1_weights[434][3] = -2;
        layer_1_weights[435][3] = 0;
        layer_1_weights[436][3] = 2;
        layer_1_weights[437][3] = 2;
        layer_1_weights[438][3] = 3;
        layer_1_weights[439][3] = 1;
        layer_1_weights[440][3] = 0;
        layer_1_weights[441][3] = 1;
        layer_1_weights[442][3] = 0;
        layer_1_weights[443][3] = 3;
        layer_1_weights[444][3] = 3;
        layer_1_weights[445][3] = 2;
        layer_1_weights[446][3] = -2;
        layer_1_weights[447][3] = -1;
        layer_1_weights[448][3] = 2;
        layer_1_weights[449][3] = -2;
        layer_1_weights[450][3] = 0;
        layer_1_weights[451][3] = -1;
        layer_1_weights[452][3] = 1;
        layer_1_weights[453][3] = 2;
        layer_1_weights[454][3] = 0;
        layer_1_weights[455][3] = 0;
        layer_1_weights[456][3] = 2;
        layer_1_weights[457][3] = 1;
        layer_1_weights[458][3] = 0;
        layer_1_weights[459][3] = -1;
        layer_1_weights[460][3] = -2;
        layer_1_weights[461][3] = -1;
        layer_1_weights[462][3] = 0;
        layer_1_weights[463][3] = 2;
        layer_1_weights[464][3] = 2;
        layer_1_weights[465][3] = 2;
        layer_1_weights[466][3] = 1;
        layer_1_weights[467][3] = 1;
        layer_1_weights[468][3] = 1;
        layer_1_weights[469][3] = 2;
        layer_1_weights[470][3] = 1;
        layer_1_weights[471][3] = 1;
        layer_1_weights[472][3] = -1;
        layer_1_weights[473][3] = 0;
        layer_1_weights[474][3] = -1;
        layer_1_weights[475][3] = -2;
        layer_1_weights[476][3] = 0;
        layer_1_weights[477][3] = -3;
        layer_1_weights[478][3] = 1;
        layer_1_weights[479][3] = 0;
        layer_1_weights[480][3] = 1;
        layer_1_weights[481][3] = 1;
        layer_1_weights[482][3] = 1;
        layer_1_weights[483][3] = 1;
        layer_1_weights[484][3] = 0;
        layer_1_weights[485][3] = 1;
        layer_1_weights[486][3] = -1;
        layer_1_weights[487][3] = -1;
        layer_1_weights[488][3] = -1;
        layer_1_weights[489][3] = 0;
        layer_1_weights[490][3] = 0;
        layer_1_weights[491][3] = 2;
        layer_1_weights[492][3] = 2;
        layer_1_weights[493][3] = 2;
        layer_1_weights[494][3] = 2;
        layer_1_weights[495][3] = 1;
        layer_1_weights[496][3] = 2;
        layer_1_weights[497][3] = 1;
        layer_1_weights[498][3] = 0;
        layer_1_weights[499][3] = 1;
        layer_1_weights[500][3] = 4;
        layer_1_weights[501][3] = 6;
        layer_1_weights[502][3] = 4;
        layer_1_weights[503][3] = -2;
        layer_1_weights[504][3] = 1;
        layer_1_weights[505][3] = 2;
        layer_1_weights[506][3] = 3;
        layer_1_weights[507][3] = -2;
        layer_1_weights[508][3] = 3;
        layer_1_weights[509][3] = 0;
        layer_1_weights[510][3] = 1;
        layer_1_weights[511][3] = 1;
        layer_1_weights[512][3] = -1;
        layer_1_weights[513][3] = -1;
        layer_1_weights[514][3] = -2;
        layer_1_weights[515][3] = -2;
        layer_1_weights[516][3] = -1;
        layer_1_weights[517][3] = 1;
        layer_1_weights[518][3] = 2;
        layer_1_weights[519][3] = 0;
        layer_1_weights[520][3] = 1;
        layer_1_weights[521][3] = 1;
        layer_1_weights[522][3] = 1;
        layer_1_weights[523][3] = 0;
        layer_1_weights[524][3] = 0;
        layer_1_weights[525][3] = 0;
        layer_1_weights[526][3] = -2;
        layer_1_weights[527][3] = 0;
        layer_1_weights[528][3] = 4;
        layer_1_weights[529][3] = 4;
        layer_1_weights[530][3] = 3;
        layer_1_weights[531][3] = -2;
        layer_1_weights[532][3] = -1;
        layer_1_weights[533][3] = 3;
        layer_1_weights[534][3] = 1;
        layer_1_weights[535][3] = 1;
        layer_1_weights[536][3] = -1;
        layer_1_weights[537][3] = -1;
        layer_1_weights[538][3] = 0;
        layer_1_weights[539][3] = -1;
        layer_1_weights[540][3] = 0;
        layer_1_weights[541][3] = -2;
        layer_1_weights[542][3] = -1;
        layer_1_weights[543][3] = -1;
        layer_1_weights[544][3] = 0;
        layer_1_weights[545][3] = 1;
        layer_1_weights[546][3] = 1;
        layer_1_weights[547][3] = 1;
        layer_1_weights[548][3] = 0;
        layer_1_weights[549][3] = -1;
        layer_1_weights[550][3] = -1;
        layer_1_weights[551][3] = 0;
        layer_1_weights[552][3] = 0;
        layer_1_weights[553][3] = -2;
        layer_1_weights[554][3] = -1;
        layer_1_weights[555][3] = -3;
        layer_1_weights[556][3] = 1;
        layer_1_weights[557][3] = 1;
        layer_1_weights[558][3] = -1;
        layer_1_weights[559][3] = -1;
        layer_1_weights[560][3] = 0;
        layer_1_weights[561][3] = 0;
        layer_1_weights[562][3] = 1;
        layer_1_weights[563][3] = -2;
        layer_1_weights[564][3] = 0;
        layer_1_weights[565][3] = -1;
        layer_1_weights[566][3] = -3;
        layer_1_weights[567][3] = -1;
        layer_1_weights[568][3] = 0;
        layer_1_weights[569][3] = 0;
        layer_1_weights[570][3] = -1;
        layer_1_weights[571][3] = 0;
        layer_1_weights[572][3] = 1;
        layer_1_weights[573][3] = 1;
        layer_1_weights[574][3] = 1;
        layer_1_weights[575][3] = -1;
        layer_1_weights[576][3] = -1;
        layer_1_weights[577][3] = -2;
        layer_1_weights[578][3] = -3;
        layer_1_weights[579][3] = 0;
        layer_1_weights[580][3] = -2;
        layer_1_weights[581][3] = -2;
        layer_1_weights[582][3] = 0;
        layer_1_weights[583][3] = -2;
        layer_1_weights[584][3] = -2;
        layer_1_weights[585][3] = -3;
        layer_1_weights[586][3] = -1;
        layer_1_weights[587][3] = 1;
        layer_1_weights[588][3] = 0;
        layer_1_weights[589][3] = -1;
        layer_1_weights[590][3] = -2;
        layer_1_weights[591][3] = -3;
        layer_1_weights[592][3] = 1;
        layer_1_weights[593][3] = -1;
        layer_1_weights[594][3] = -3;
        layer_1_weights[595][3] = -1;
        layer_1_weights[596][3] = 0;
        layer_1_weights[597][3] = -1;
        layer_1_weights[598][3] = 0;
        layer_1_weights[599][3] = 1;
        layer_1_weights[600][3] = -1;
        layer_1_weights[601][3] = -1;
        layer_1_weights[602][3] = 0;
        layer_1_weights[603][3] = 0;
        layer_1_weights[604][3] = -1;
        layer_1_weights[605][3] = -1;
        layer_1_weights[606][3] = -1;
        layer_1_weights[607][3] = -2;
        layer_1_weights[608][3] = -2;
        layer_1_weights[609][3] = 0;
        layer_1_weights[610][3] = 2;
        layer_1_weights[611][3] = -1;
        layer_1_weights[612][3] = 0;
        layer_1_weights[613][3] = -1;
        layer_1_weights[614][3] = 1;
        layer_1_weights[615][3] = 1;
        layer_1_weights[616][3] = -1;
        layer_1_weights[617][3] = 0;
        layer_1_weights[618][3] = -4;
        layer_1_weights[619][3] = -5;
        layer_1_weights[620][3] = -2;
        layer_1_weights[621][3] = -1;
        layer_1_weights[622][3] = -1;
        layer_1_weights[623][3] = 0;
        layer_1_weights[624][3] = -1;
        layer_1_weights[625][3] = 1;
        layer_1_weights[626][3] = -1;
        layer_1_weights[627][3] = 1;
        layer_1_weights[628][3] = 1;
        layer_1_weights[629][3] = 1;
        layer_1_weights[630][3] = -1;
        layer_1_weights[631][3] = 0;
        layer_1_weights[632][3] = 1;
        layer_1_weights[633][3] = 0;
        layer_1_weights[634][3] = -1;
        layer_1_weights[635][3] = -1;
        layer_1_weights[636][3] = 1;
        layer_1_weights[637][3] = -2;
        layer_1_weights[638][3] = 1;
        layer_1_weights[639][3] = 0;
        layer_1_weights[640][3] = 1;
        layer_1_weights[641][3] = 1;
        layer_1_weights[642][3] = 1;
        layer_1_weights[643][3] = 1;
        layer_1_weights[644][3] = 1;
        layer_1_weights[645][3] = -1;
        layer_1_weights[646][3] = -3;
        layer_1_weights[647][3] = -3;
        layer_1_weights[648][3] = -2;
        layer_1_weights[649][3] = -1;
        layer_1_weights[650][3] = 0;
        layer_1_weights[651][3] = 0;
        layer_1_weights[652][3] = 1;
        layer_1_weights[653][3] = 1;
        layer_1_weights[654][3] = 0;
        layer_1_weights[655][3] = 0;
        layer_1_weights[656][3] = 1;
        layer_1_weights[657][3] = 0;
        layer_1_weights[658][3] = -1;
        layer_1_weights[659][3] = -1;
        layer_1_weights[660][3] = 1;
        layer_1_weights[661][3] = 0;
        layer_1_weights[662][3] = -2;
        layer_1_weights[663][3] = -1;
        layer_1_weights[664][3] = 0;
        layer_1_weights[665][3] = -1;
        layer_1_weights[666][3] = 0;
        layer_1_weights[667][3] = -2;
        layer_1_weights[668][3] = 1;
        layer_1_weights[669][3] = 2;
        layer_1_weights[670][3] = 2;
        layer_1_weights[671][3] = 0;
        layer_1_weights[672][3] = 0;
        layer_1_weights[673][3] = 0;
        layer_1_weights[674][3] = 2;
        layer_1_weights[675][3] = 1;
        layer_1_weights[676][3] = -1;
        layer_1_weights[677][3] = 0;
        layer_1_weights[678][3] = -2;
        layer_1_weights[679][3] = -1;
        layer_1_weights[680][3] = 0;
        layer_1_weights[681][3] = 0;
        layer_1_weights[682][3] = -1;
        layer_1_weights[683][3] = 0;
        layer_1_weights[684][3] = 0;
        layer_1_weights[685][3] = -1;
        layer_1_weights[686][3] = 1;
        layer_1_weights[687][3] = 1;
        layer_1_weights[688][3] = 2;
        layer_1_weights[689][3] = 0;
        layer_1_weights[690][3] = 1;
        layer_1_weights[691][3] = 0;
        layer_1_weights[692][3] = 1;
        layer_1_weights[693][3] = 2;
        layer_1_weights[694][3] = 2;
        layer_1_weights[695][3] = -2;
        layer_1_weights[696][3] = 1;
        layer_1_weights[697][3] = 0;
        layer_1_weights[698][3] = 1;
        layer_1_weights[699][3] = 0;
        layer_1_weights[700][3] = -1;
        layer_1_weights[701][3] = 0;
        layer_1_weights[702][3] = -3;
        layer_1_weights[703][3] = 2;
        layer_1_weights[704][3] = -1;
        layer_1_weights[705][3] = 0;
        layer_1_weights[706][3] = -1;
        layer_1_weights[707][3] = -1;
        layer_1_weights[708][3] = -2;
        layer_1_weights[709][3] = -2;
        layer_1_weights[710][3] = -1;
        layer_1_weights[711][3] = 0;
        layer_1_weights[712][3] = -1;
        layer_1_weights[713][3] = 0;
        layer_1_weights[714][3] = 1;
        layer_1_weights[715][3] = 2;
        layer_1_weights[716][3] = 2;
        layer_1_weights[717][3] = 2;
        layer_1_weights[718][3] = 2;
        layer_1_weights[719][3] = 0;
        layer_1_weights[720][3] = 0;
        layer_1_weights[721][3] = 1;
        layer_1_weights[722][3] = 0;
        layer_1_weights[723][3] = 0;
        layer_1_weights[724][3] = 1;
        layer_1_weights[725][3] = -2;
        layer_1_weights[726][3] = 0;
        layer_1_weights[727][3] = 0;
        layer_1_weights[728][3] = 0;
        layer_1_weights[729][3] = -1;
        layer_1_weights[730][3] = 0;
        layer_1_weights[731][3] = 0;
        layer_1_weights[732][3] = -1;
        layer_1_weights[733][3] = -3;
        layer_1_weights[734][3] = -3;
        layer_1_weights[735][3] = -3;
        layer_1_weights[736][3] = -3;
        layer_1_weights[737][3] = -1;
        layer_1_weights[738][3] = -2;
        layer_1_weights[739][3] = -1;
        layer_1_weights[740][3] = -1;
        layer_1_weights[741][3] = 2;
        layer_1_weights[742][3] = 0;
        layer_1_weights[743][3] = 0;
        layer_1_weights[744][3] = 1;
        layer_1_weights[745][3] = 1;
        layer_1_weights[746][3] = 1;
        layer_1_weights[747][3] = 2;
        layer_1_weights[748][3] = 0;
        layer_1_weights[749][3] = 0;
        layer_1_weights[750][3] = 1;
        layer_1_weights[751][3] = -1;
        layer_1_weights[752][3] = 0;
        layer_1_weights[753][3] = 2;
        layer_1_weights[754][3] = 0;
        layer_1_weights[755][3] = -1;
        layer_1_weights[756][3] = 0;
        layer_1_weights[757][3] = 0;
        layer_1_weights[758][3] = 0;
        layer_1_weights[759][3] = 0;
        layer_1_weights[760][3] = 3;
        layer_1_weights[761][3] = 4;
        layer_1_weights[762][3] = -2;
        layer_1_weights[763][3] = -1;
        layer_1_weights[764][3] = -1;
        layer_1_weights[765][3] = -2;
        layer_1_weights[766][3] = 1;
        layer_1_weights[767][3] = 0;
        layer_1_weights[768][3] = 1;
        layer_1_weights[769][3] = 3;
        layer_1_weights[770][3] = -1;
        layer_1_weights[771][3] = 0;
        layer_1_weights[772][3] = 0;
        layer_1_weights[773][3] = 2;
        layer_1_weights[774][3] = -1;
        layer_1_weights[775][3] = 2;
        layer_1_weights[776][3] = -1;
        layer_1_weights[777][3] = 3;
        layer_1_weights[778][3] = 1;
        layer_1_weights[779][3] = 3;
        layer_1_weights[780][3] = 0;
        layer_1_weights[781][3] = 0;
        layer_1_weights[782][3] = -1;
        layer_1_weights[783][3] = 0;
        layer_1_weights[0][4] = 0;
        layer_1_weights[1][4] = 1;
        layer_1_weights[2][4] = 0;
        layer_1_weights[3][4] = 0;
        layer_1_weights[4][4] = 0;
        layer_1_weights[5][4] = 1;
        layer_1_weights[6][4] = 0;
        layer_1_weights[7][4] = 0;
        layer_1_weights[8][4] = -1;
        layer_1_weights[9][4] = 0;
        layer_1_weights[10][4] = 0;
        layer_1_weights[11][4] = 0;
        layer_1_weights[12][4] = -1;
        layer_1_weights[13][4] = -1;
        layer_1_weights[14][4] = 0;
        layer_1_weights[15][4] = 1;
        layer_1_weights[16][4] = -1;
        layer_1_weights[17][4] = 1;
        layer_1_weights[18][4] = 0;
        layer_1_weights[19][4] = 0;
        layer_1_weights[20][4] = 0;
        layer_1_weights[21][4] = 0;
        layer_1_weights[22][4] = 0;
        layer_1_weights[23][4] = 0;
        layer_1_weights[24][4] = 0;
        layer_1_weights[25][4] = 0;
        layer_1_weights[26][4] = 0;
        layer_1_weights[27][4] = 0;
        layer_1_weights[28][4] = -1;
        layer_1_weights[29][4] = 1;
        layer_1_weights[30][4] = 1;
        layer_1_weights[31][4] = 0;
        layer_1_weights[32][4] = 1;
        layer_1_weights[33][4] = -1;
        layer_1_weights[34][4] = -3;
        layer_1_weights[35][4] = -2;
        layer_1_weights[36][4] = -3;
        layer_1_weights[37][4] = -3;
        layer_1_weights[38][4] = -4;
        layer_1_weights[39][4] = -4;
        layer_1_weights[40][4] = -4;
        layer_1_weights[41][4] = -4;
        layer_1_weights[42][4] = -2;
        layer_1_weights[43][4] = -2;
        layer_1_weights[44][4] = 0;
        layer_1_weights[45][4] = -2;
        layer_1_weights[46][4] = -2;
        layer_1_weights[47][4] = -3;
        layer_1_weights[48][4] = -2;
        layer_1_weights[49][4] = -1;
        layer_1_weights[50][4] = -2;
        layer_1_weights[51][4] = -1;
        layer_1_weights[52][4] = -1;
        layer_1_weights[53][4] = 0;
        layer_1_weights[54][4] = 0;
        layer_1_weights[55][4] = 0;
        layer_1_weights[56][4] = 0;
        layer_1_weights[57][4] = 0;
        layer_1_weights[58][4] = 1;
        layer_1_weights[59][4] = -1;
        layer_1_weights[60][4] = -1;
        layer_1_weights[61][4] = 0;
        layer_1_weights[62][4] = -4;
        layer_1_weights[63][4] = -6;
        layer_1_weights[64][4] = -1;
        layer_1_weights[65][4] = 0;
        layer_1_weights[66][4] = -1;
        layer_1_weights[67][4] = 0;
        layer_1_weights[68][4] = -2;
        layer_1_weights[69][4] = -5;
        layer_1_weights[70][4] = -2;
        layer_1_weights[71][4] = -5;
        layer_1_weights[72][4] = -2;
        layer_1_weights[73][4] = 0;
        layer_1_weights[74][4] = -1;
        layer_1_weights[75][4] = -2;
        layer_1_weights[76][4] = -4;
        layer_1_weights[77][4] = -2;
        layer_1_weights[78][4] = -2;
        layer_1_weights[79][4] = 1;
        layer_1_weights[80][4] = 3;
        layer_1_weights[81][4] = 0;
        layer_1_weights[82][4] = 0;
        layer_1_weights[83][4] = 0;
        layer_1_weights[84][4] = 0;
        layer_1_weights[85][4] = 0;
        layer_1_weights[86][4] = -1;
        layer_1_weights[87][4] = -2;
        layer_1_weights[88][4] = -1;
        layer_1_weights[89][4] = 2;
        layer_1_weights[90][4] = 4;
        layer_1_weights[91][4] = 3;
        layer_1_weights[92][4] = -1;
        layer_1_weights[93][4] = -4;
        layer_1_weights[94][4] = -3;
        layer_1_weights[95][4] = -4;
        layer_1_weights[96][4] = -3;
        layer_1_weights[97][4] = -6;
        layer_1_weights[98][4] = -6;
        layer_1_weights[99][4] = -5;
        layer_1_weights[100][4] = -5;
        layer_1_weights[101][4] = -3;
        layer_1_weights[102][4] = -3;
        layer_1_weights[103][4] = -3;
        layer_1_weights[104][4] = -1;
        layer_1_weights[105][4] = -2;
        layer_1_weights[106][4] = 1;
        layer_1_weights[107][4] = 2;
        layer_1_weights[108][4] = 2;
        layer_1_weights[109][4] = 2;
        layer_1_weights[110][4] = 1;
        layer_1_weights[111][4] = 0;
        layer_1_weights[112][4] = 0;
        layer_1_weights[113][4] = 2;
        layer_1_weights[114][4] = 0;
        layer_1_weights[115][4] = -1;
        layer_1_weights[116][4] = 0;
        layer_1_weights[117][4] = 3;
        layer_1_weights[118][4] = 2;
        layer_1_weights[119][4] = 1;
        layer_1_weights[120][4] = -1;
        layer_1_weights[121][4] = -1;
        layer_1_weights[122][4] = 0;
        layer_1_weights[123][4] = 1;
        layer_1_weights[124][4] = 1;
        layer_1_weights[125][4] = -1;
        layer_1_weights[126][4] = -1;
        layer_1_weights[127][4] = -2;
        layer_1_weights[128][4] = -4;
        layer_1_weights[129][4] = -3;
        layer_1_weights[130][4] = -1;
        layer_1_weights[131][4] = -2;
        layer_1_weights[132][4] = -4;
        layer_1_weights[133][4] = -3;
        layer_1_weights[134][4] = -1;
        layer_1_weights[135][4] = -1;
        layer_1_weights[136][4] = 2;
        layer_1_weights[137][4] = 5;
        layer_1_weights[138][4] = 2;
        layer_1_weights[139][4] = 1;
        layer_1_weights[140][4] = 1;
        layer_1_weights[141][4] = 0;
        layer_1_weights[142][4] = -2;
        layer_1_weights[143][4] = 1;
        layer_1_weights[144][4] = -1;
        layer_1_weights[145][4] = 2;
        layer_1_weights[146][4] = 1;
        layer_1_weights[147][4] = 1;
        layer_1_weights[148][4] = 1;
        layer_1_weights[149][4] = 1;
        layer_1_weights[150][4] = 1;
        layer_1_weights[151][4] = 0;
        layer_1_weights[152][4] = 1;
        layer_1_weights[153][4] = 2;
        layer_1_weights[154][4] = -1;
        layer_1_weights[155][4] = -1;
        layer_1_weights[156][4] = 0;
        layer_1_weights[157][4] = -2;
        layer_1_weights[158][4] = -3;
        layer_1_weights[159][4] = -2;
        layer_1_weights[160][4] = -1;
        layer_1_weights[161][4] = -1;
        layer_1_weights[162][4] = -1;
        layer_1_weights[163][4] = -1;
        layer_1_weights[164][4] = 2;
        layer_1_weights[165][4] = 5;
        layer_1_weights[166][4] = -1;
        layer_1_weights[167][4] = 1;
        layer_1_weights[168][4] = 0;
        layer_1_weights[169][4] = -1;
        layer_1_weights[170][4] = 2;
        layer_1_weights[171][4] = 6;
        layer_1_weights[172][4] = 2;
        layer_1_weights[173][4] = 2;
        layer_1_weights[174][4] = 2;
        layer_1_weights[175][4] = 1;
        layer_1_weights[176][4] = 1;
        layer_1_weights[177][4] = 1;
        layer_1_weights[178][4] = 1;
        layer_1_weights[179][4] = 2;
        layer_1_weights[180][4] = 2;
        layer_1_weights[181][4] = 2;
        layer_1_weights[182][4] = 1;
        layer_1_weights[183][4] = 1;
        layer_1_weights[184][4] = 2;
        layer_1_weights[185][4] = 0;
        layer_1_weights[186][4] = -2;
        layer_1_weights[187][4] = -3;
        layer_1_weights[188][4] = -2;
        layer_1_weights[189][4] = 0;
        layer_1_weights[190][4] = -2;
        layer_1_weights[191][4] = -2;
        layer_1_weights[192][4] = 1;
        layer_1_weights[193][4] = 5;
        layer_1_weights[194][4] = 2;
        layer_1_weights[195][4] = 3;
        layer_1_weights[196][4] = 0;
        layer_1_weights[197][4] = 1;
        layer_1_weights[198][4] = 2;
        layer_1_weights[199][4] = 5;
        layer_1_weights[200][4] = 4;
        layer_1_weights[201][4] = 2;
        layer_1_weights[202][4] = 3;
        layer_1_weights[203][4] = 0;
        layer_1_weights[204][4] = 1;
        layer_1_weights[205][4] = 1;
        layer_1_weights[206][4] = 1;
        layer_1_weights[207][4] = 2;
        layer_1_weights[208][4] = 1;
        layer_1_weights[209][4] = 2;
        layer_1_weights[210][4] = 2;
        layer_1_weights[211][4] = 1;
        layer_1_weights[212][4] = 2;
        layer_1_weights[213][4] = 0;
        layer_1_weights[214][4] = -2;
        layer_1_weights[215][4] = -3;
        layer_1_weights[216][4] = -1;
        layer_1_weights[217][4] = -1;
        layer_1_weights[218][4] = -1;
        layer_1_weights[219][4] = 0;
        layer_1_weights[220][4] = 2;
        layer_1_weights[221][4] = 5;
        layer_1_weights[222][4] = 2;
        layer_1_weights[223][4] = 3;
        layer_1_weights[224][4] = -3;
        layer_1_weights[225][4] = 2;
        layer_1_weights[226][4] = 1;
        layer_1_weights[227][4] = 3;
        layer_1_weights[228][4] = 6;
        layer_1_weights[229][4] = 0;
        layer_1_weights[230][4] = 1;
        layer_1_weights[231][4] = 1;
        layer_1_weights[232][4] = 2;
        layer_1_weights[233][4] = 2;
        layer_1_weights[234][4] = 1;
        layer_1_weights[235][4] = 0;
        layer_1_weights[236][4] = 1;
        layer_1_weights[237][4] = 2;
        layer_1_weights[238][4] = 4;
        layer_1_weights[239][4] = 3;
        layer_1_weights[240][4] = 1;
        layer_1_weights[241][4] = 0;
        layer_1_weights[242][4] = 0;
        layer_1_weights[243][4] = -3;
        layer_1_weights[244][4] = -2;
        layer_1_weights[245][4] = -1;
        layer_1_weights[246][4] = -2;
        layer_1_weights[247][4] = -2;
        layer_1_weights[248][4] = 0;
        layer_1_weights[249][4] = 1;
        layer_1_weights[250][4] = 4;
        layer_1_weights[251][4] = -1;
        layer_1_weights[252][4] = 1;
        layer_1_weights[253][4] = 1;
        layer_1_weights[254][4] = 3;
        layer_1_weights[255][4] = 5;
        layer_1_weights[256][4] = 2;
        layer_1_weights[257][4] = 0;
        layer_1_weights[258][4] = 1;
        layer_1_weights[259][4] = 1;
        layer_1_weights[260][4] = 1;
        layer_1_weights[261][4] = 1;
        layer_1_weights[262][4] = 1;
        layer_1_weights[263][4] = 2;
        layer_1_weights[264][4] = 2;
        layer_1_weights[265][4] = 2;
        layer_1_weights[266][4] = 3;
        layer_1_weights[267][4] = 3;
        layer_1_weights[268][4] = 1;
        layer_1_weights[269][4] = 1;
        layer_1_weights[270][4] = 0;
        layer_1_weights[271][4] = -1;
        layer_1_weights[272][4] = -1;
        layer_1_weights[273][4] = -2;
        layer_1_weights[274][4] = -2;
        layer_1_weights[275][4] = -2;
        layer_1_weights[276][4] = -1;
        layer_1_weights[277][4] = 1;
        layer_1_weights[278][4] = 4;
        layer_1_weights[279][4] = 3;
        layer_1_weights[280][4] = 1;
        layer_1_weights[281][4] = -1;
        layer_1_weights[282][4] = 4;
        layer_1_weights[283][4] = 8;
        layer_1_weights[284][4] = 0;
        layer_1_weights[285][4] = 1;
        layer_1_weights[286][4] = 1;
        layer_1_weights[287][4] = -1;
        layer_1_weights[288][4] = -1;
        layer_1_weights[289][4] = 0;
        layer_1_weights[290][4] = -1;
        layer_1_weights[291][4] = -2;
        layer_1_weights[292][4] = -1;
        layer_1_weights[293][4] = -1;
        layer_1_weights[294][4] = -1;
        layer_1_weights[295][4] = 0;
        layer_1_weights[296][4] = 1;
        layer_1_weights[297][4] = 2;
        layer_1_weights[298][4] = 2;
        layer_1_weights[299][4] = 1;
        layer_1_weights[300][4] = 1;
        layer_1_weights[301][4] = -2;
        layer_1_weights[302][4] = -3;
        layer_1_weights[303][4] = -1;
        layer_1_weights[304][4] = -3;
        layer_1_weights[305][4] = 2;
        layer_1_weights[306][4] = -1;
        layer_1_weights[307][4] = 2;
        layer_1_weights[308][4] = 0;
        layer_1_weights[309][4] = -2;
        layer_1_weights[310][4] = 3;
        layer_1_weights[311][4] = 5;
        layer_1_weights[312][4] = -2;
        layer_1_weights[313][4] = 0;
        layer_1_weights[314][4] = -1;
        layer_1_weights[315][4] = -1;
        layer_1_weights[316][4] = -1;
        layer_1_weights[317][4] = 0;
        layer_1_weights[318][4] = -1;
        layer_1_weights[319][4] = -1;
        layer_1_weights[320][4] = -1;
        layer_1_weights[321][4] = -1;
        layer_1_weights[322][4] = -1;
        layer_1_weights[323][4] = 1;
        layer_1_weights[324][4] = 2;
        layer_1_weights[325][4] = 3;
        layer_1_weights[326][4] = 3;
        layer_1_weights[327][4] = 2;
        layer_1_weights[328][4] = 1;
        layer_1_weights[329][4] = 0;
        layer_1_weights[330][4] = -2;
        layer_1_weights[331][4] = -2;
        layer_1_weights[332][4] = -3;
        layer_1_weights[333][4] = -3;
        layer_1_weights[334][4] = 0;
        layer_1_weights[335][4] = 1;
        layer_1_weights[336][4] = 0;
        layer_1_weights[337][4] = 1;
        layer_1_weights[338][4] = 4;
        layer_1_weights[339][4] = 3;
        layer_1_weights[340][4] = -3;
        layer_1_weights[341][4] = -3;
        layer_1_weights[342][4] = -3;
        layer_1_weights[343][4] = -2;
        layer_1_weights[344][4] = -2;
        layer_1_weights[345][4] = -1;
        layer_1_weights[346][4] = -1;
        layer_1_weights[347][4] = -2;
        layer_1_weights[348][4] = -2;
        layer_1_weights[349][4] = -1;
        layer_1_weights[350][4] = 0;
        layer_1_weights[351][4] = 1;
        layer_1_weights[352][4] = 2;
        layer_1_weights[353][4] = 2;
        layer_1_weights[354][4] = 5;
        layer_1_weights[355][4] = 3;
        layer_1_weights[356][4] = -1;
        layer_1_weights[357][4] = -2;
        layer_1_weights[358][4] = -2;
        layer_1_weights[359][4] = -6;
        layer_1_weights[360][4] = -3;
        layer_1_weights[361][4] = -2;
        layer_1_weights[362][4] = -1;
        layer_1_weights[363][4] = -1;
        layer_1_weights[364][4] = 0;
        layer_1_weights[365][4] = -1;
        layer_1_weights[366][4] = 0;
        layer_1_weights[367][4] = 1;
        layer_1_weights[368][4] = -3;
        layer_1_weights[369][4] = -4;
        layer_1_weights[370][4] = -2;
        layer_1_weights[371][4] = -1;
        layer_1_weights[372][4] = -1;
        layer_1_weights[373][4] = 0;
        layer_1_weights[374][4] = 1;
        layer_1_weights[375][4] = 1;
        layer_1_weights[376][4] = 1;
        layer_1_weights[377][4] = 0;
        layer_1_weights[378][4] = 2;
        layer_1_weights[379][4] = 2;
        layer_1_weights[380][4] = 2;
        layer_1_weights[381][4] = 2;
        layer_1_weights[382][4] = 2;
        layer_1_weights[383][4] = 1;
        layer_1_weights[384][4] = -2;
        layer_1_weights[385][4] = -3;
        layer_1_weights[386][4] = -4;
        layer_1_weights[387][4] = -1;
        layer_1_weights[388][4] = -2;
        layer_1_weights[389][4] = 3;
        layer_1_weights[390][4] = 4;
        layer_1_weights[391][4] = 0;
        layer_1_weights[392][4] = -2;
        layer_1_weights[393][4] = 1;
        layer_1_weights[394][4] = 4;
        layer_1_weights[395][4] = 2;
        layer_1_weights[396][4] = -2;
        layer_1_weights[397][4] = -4;
        layer_1_weights[398][4] = -1;
        layer_1_weights[399][4] = 0;
        layer_1_weights[400][4] = -1;
        layer_1_weights[401][4] = 0;
        layer_1_weights[402][4] = -1;
        layer_1_weights[403][4] = 1;
        layer_1_weights[404][4] = 0;
        layer_1_weights[405][4] = 1;
        layer_1_weights[406][4] = 1;
        layer_1_weights[407][4] = 3;
        layer_1_weights[408][4] = 3;
        layer_1_weights[409][4] = 2;
        layer_1_weights[410][4] = 3;
        layer_1_weights[411][4] = 1;
        layer_1_weights[412][4] = -2;
        layer_1_weights[413][4] = -2;
        layer_1_weights[414][4] = -2;
        layer_1_weights[415][4] = -1;
        layer_1_weights[416][4] = -1;
        layer_1_weights[417][4] = 2;
        layer_1_weights[418][4] = 5;
        layer_1_weights[419][4] = 0;
        layer_1_weights[420][4] = -2;
        layer_1_weights[421][4] = 2;
        layer_1_weights[422][4] = 0;
        layer_1_weights[423][4] = 3;
        layer_1_weights[424][4] = -1;
        layer_1_weights[425][4] = -2;
        layer_1_weights[426][4] = 0;
        layer_1_weights[427][4] = 0;
        layer_1_weights[428][4] = -2;
        layer_1_weights[429][4] = -1;
        layer_1_weights[430][4] = 0;
        layer_1_weights[431][4] = 0;
        layer_1_weights[432][4] = 0;
        layer_1_weights[433][4] = 0;
        layer_1_weights[434][4] = 1;
        layer_1_weights[435][4] = 3;
        layer_1_weights[436][4] = 3;
        layer_1_weights[437][4] = 2;
        layer_1_weights[438][4] = -1;
        layer_1_weights[439][4] = -2;
        layer_1_weights[440][4] = -1;
        layer_1_weights[441][4] = -1;
        layer_1_weights[442][4] = 1;
        layer_1_weights[443][4] = -1;
        layer_1_weights[444][4] = 3;
        layer_1_weights[445][4] = 0;
        layer_1_weights[446][4] = 9;
        layer_1_weights[447][4] = 3;
        layer_1_weights[448][4] = 3;
        layer_1_weights[449][4] = 2;
        layer_1_weights[450][4] = 1;
        layer_1_weights[451][4] = 4;
        layer_1_weights[452][4] = 0;
        layer_1_weights[453][4] = -3;
        layer_1_weights[454][4] = -2;
        layer_1_weights[455][4] = -1;
        layer_1_weights[456][4] = -2;
        layer_1_weights[457][4] = -1;
        layer_1_weights[458][4] = -1;
        layer_1_weights[459][4] = 1;
        layer_1_weights[460][4] = 1;
        layer_1_weights[461][4] = 1;
        layer_1_weights[462][4] = 1;
        layer_1_weights[463][4] = 2;
        layer_1_weights[464][4] = 2;
        layer_1_weights[465][4] = 2;
        layer_1_weights[466][4] = 0;
        layer_1_weights[467][4] = -1;
        layer_1_weights[468][4] = 0;
        layer_1_weights[469][4] = 0;
        layer_1_weights[470][4] = 3;
        layer_1_weights[471][4] = 1;
        layer_1_weights[472][4] = 4;
        layer_1_weights[473][4] = 1;
        layer_1_weights[474][4] = 7;
        layer_1_weights[475][4] = 4;
        layer_1_weights[476][4] = 0;
        layer_1_weights[477][4] = 2;
        layer_1_weights[478][4] = 2;
        layer_1_weights[479][4] = 0;
        layer_1_weights[480][4] = 0;
        layer_1_weights[481][4] = -2;
        layer_1_weights[482][4] = -2;
        layer_1_weights[483][4] = 0;
        layer_1_weights[484][4] = 0;
        layer_1_weights[485][4] = -1;
        layer_1_weights[486][4] = -1;
        layer_1_weights[487][4] = 0;
        layer_1_weights[488][4] = -1;
        layer_1_weights[489][4] = 1;
        layer_1_weights[490][4] = 0;
        layer_1_weights[491][4] = 1;
        layer_1_weights[492][4] = 0;
        layer_1_weights[493][4] = -1;
        layer_1_weights[494][4] = -1;
        layer_1_weights[495][4] = -3;
        layer_1_weights[496][4] = -1;
        layer_1_weights[497][4] = -2;
        layer_1_weights[498][4] = 1;
        layer_1_weights[499][4] = 0;
        layer_1_weights[500][4] = -2;
        layer_1_weights[501][4] = 5;
        layer_1_weights[502][4] = 2;
        layer_1_weights[503][4] = 2;
        layer_1_weights[504][4] = 3;
        layer_1_weights[505][4] = 2;
        layer_1_weights[506][4] = 4;
        layer_1_weights[507][4] = 3;
        layer_1_weights[508][4] = 1;
        layer_1_weights[509][4] = 0;
        layer_1_weights[510][4] = 2;
        layer_1_weights[511][4] = -1;
        layer_1_weights[512][4] = 0;
        layer_1_weights[513][4] = -1;
        layer_1_weights[514][4] = -1;
        layer_1_weights[515][4] = 1;
        layer_1_weights[516][4] = 0;
        layer_1_weights[517][4] = -1;
        layer_1_weights[518][4] = 0;
        layer_1_weights[519][4] = 0;
        layer_1_weights[520][4] = -2;
        layer_1_weights[521][4] = -2;
        layer_1_weights[522][4] = 0;
        layer_1_weights[523][4] = -1;
        layer_1_weights[524][4] = -1;
        layer_1_weights[525][4] = 1;
        layer_1_weights[526][4] = 0;
        layer_1_weights[527][4] = -1;
        layer_1_weights[528][4] = -2;
        layer_1_weights[529][4] = -1;
        layer_1_weights[530][4] = 1;
        layer_1_weights[531][4] = 1;
        layer_1_weights[532][4] = 0;
        layer_1_weights[533][4] = 2;
        layer_1_weights[534][4] = 2;
        layer_1_weights[535][4] = 5;
        layer_1_weights[536][4] = 2;
        layer_1_weights[537][4] = 0;
        layer_1_weights[538][4] = 0;
        layer_1_weights[539][4] = -1;
        layer_1_weights[540][4] = -2;
        layer_1_weights[541][4] = -1;
        layer_1_weights[542][4] = -2;
        layer_1_weights[543][4] = -1;
        layer_1_weights[544][4] = -1;
        layer_1_weights[545][4] = 0;
        layer_1_weights[546][4] = 0;
        layer_1_weights[547][4] = -1;
        layer_1_weights[548][4] = -2;
        layer_1_weights[549][4] = -2;
        layer_1_weights[550][4] = -2;
        layer_1_weights[551][4] = -1;
        layer_1_weights[552][4] = -1;
        layer_1_weights[553][4] = 0;
        layer_1_weights[554][4] = -1;
        layer_1_weights[555][4] = -1;
        layer_1_weights[556][4] = -2;
        layer_1_weights[557][4] = -4;
        layer_1_weights[558][4] = 0;
        layer_1_weights[559][4] = -3;
        layer_1_weights[560][4] = 0;
        layer_1_weights[561][4] = -1;
        layer_1_weights[562][4] = 2;
        layer_1_weights[563][4] = 4;
        layer_1_weights[564][4] = 0;
        layer_1_weights[565][4] = 1;
        layer_1_weights[566][4] = 0;
        layer_1_weights[567][4] = 0;
        layer_1_weights[568][4] = -1;
        layer_1_weights[569][4] = -1;
        layer_1_weights[570][4] = -1;
        layer_1_weights[571][4] = -2;
        layer_1_weights[572][4] = 0;
        layer_1_weights[573][4] = -1;
        layer_1_weights[574][4] = -1;
        layer_1_weights[575][4] = -1;
        layer_1_weights[576][4] = -1;
        layer_1_weights[577][4] = -1;
        layer_1_weights[578][4] = -1;
        layer_1_weights[579][4] = -1;
        layer_1_weights[580][4] = 0;
        layer_1_weights[581][4] = 0;
        layer_1_weights[582][4] = -1;
        layer_1_weights[583][4] = -2;
        layer_1_weights[584][4] = -2;
        layer_1_weights[585][4] = -2;
        layer_1_weights[586][4] = -1;
        layer_1_weights[587][4] = -2;
        layer_1_weights[588][4] = 0;
        layer_1_weights[589][4] = 4;
        layer_1_weights[590][4] = 6;
        layer_1_weights[591][4] = 1;
        layer_1_weights[592][4] = -1;
        layer_1_weights[593][4] = -1;
        layer_1_weights[594][4] = -1;
        layer_1_weights[595][4] = -2;
        layer_1_weights[596][4] = 1;
        layer_1_weights[597][4] = -1;
        layer_1_weights[598][4] = 0;
        layer_1_weights[599][4] = -1;
        layer_1_weights[600][4] = 0;
        layer_1_weights[601][4] = 0;
        layer_1_weights[602][4] = 1;
        layer_1_weights[603][4] = 0;
        layer_1_weights[604][4] = 1;
        layer_1_weights[605][4] = -1;
        layer_1_weights[606][4] = -1;
        layer_1_weights[607][4] = -1;
        layer_1_weights[608][4] = -1;
        layer_1_weights[609][4] = -2;
        layer_1_weights[610][4] = -4;
        layer_1_weights[611][4] = -1;
        layer_1_weights[612][4] = -1;
        layer_1_weights[613][4] = -2;
        layer_1_weights[614][4] = -2;
        layer_1_weights[615][4] = 0;
        layer_1_weights[616][4] = 0;
        layer_1_weights[617][4] = 1;
        layer_1_weights[618][4] = 3;
        layer_1_weights[619][4] = 1;
        layer_1_weights[620][4] = -2;
        layer_1_weights[621][4] = -1;
        layer_1_weights[622][4] = -1;
        layer_1_weights[623][4] = 0;
        layer_1_weights[624][4] = -1;
        layer_1_weights[625][4] = -1;
        layer_1_weights[626][4] = 1;
        layer_1_weights[627][4] = -1;
        layer_1_weights[628][4] = 0;
        layer_1_weights[629][4] = 0;
        layer_1_weights[630][4] = 1;
        layer_1_weights[631][4] = 1;
        layer_1_weights[632][4] = 1;
        layer_1_weights[633][4] = -2;
        layer_1_weights[634][4] = 0;
        layer_1_weights[635][4] = -1;
        layer_1_weights[636][4] = -1;
        layer_1_weights[637][4] = -1;
        layer_1_weights[638][4] = -3;
        layer_1_weights[639][4] = -4;
        layer_1_weights[640][4] = -2;
        layer_1_weights[641][4] = -3;
        layer_1_weights[642][4] = -3;
        layer_1_weights[643][4] = 0;
        layer_1_weights[644][4] = 0;
        layer_1_weights[645][4] = 0;
        layer_1_weights[646][4] = 1;
        layer_1_weights[647][4] = -1;
        layer_1_weights[648][4] = -2;
        layer_1_weights[649][4] = -1;
        layer_1_weights[650][4] = 1;
        layer_1_weights[651][4] = 1;
        layer_1_weights[652][4] = -1;
        layer_1_weights[653][4] = 1;
        layer_1_weights[654][4] = 1;
        layer_1_weights[655][4] = 0;
        layer_1_weights[656][4] = 0;
        layer_1_weights[657][4] = -1;
        layer_1_weights[658][4] = 0;
        layer_1_weights[659][4] = 0;
        layer_1_weights[660][4] = 0;
        layer_1_weights[661][4] = -1;
        layer_1_weights[662][4] = 0;
        layer_1_weights[663][4] = 1;
        layer_1_weights[664][4] = -2;
        layer_1_weights[665][4] = 0;
        layer_1_weights[666][4] = 0;
        layer_1_weights[667][4] = -1;
        layer_1_weights[668][4] = 2;
        layer_1_weights[669][4] = -2;
        layer_1_weights[670][4] = -3;
        layer_1_weights[671][4] = 0;
        layer_1_weights[672][4] = -1;
        layer_1_weights[673][4] = 0;
        layer_1_weights[674][4] = 3;
        layer_1_weights[675][4] = 1;
        layer_1_weights[676][4] = 2;
        layer_1_weights[677][4] = 2;
        layer_1_weights[678][4] = 2;
        layer_1_weights[679][4] = 1;
        layer_1_weights[680][4] = 0;
        layer_1_weights[681][4] = -1;
        layer_1_weights[682][4] = -2;
        layer_1_weights[683][4] = 0;
        layer_1_weights[684][4] = -2;
        layer_1_weights[685][4] = -1;
        layer_1_weights[686][4] = 0;
        layer_1_weights[687][4] = -1;
        layer_1_weights[688][4] = 0;
        layer_1_weights[689][4] = 1;
        layer_1_weights[690][4] = 0;
        layer_1_weights[691][4] = 1;
        layer_1_weights[692][4] = -1;
        layer_1_weights[693][4] = 0;
        layer_1_weights[694][4] = -1;
        layer_1_weights[695][4] = 1;
        layer_1_weights[696][4] = -1;
        layer_1_weights[697][4] = 0;
        layer_1_weights[698][4] = -1;
        layer_1_weights[699][4] = 1;
        layer_1_weights[700][4] = -1;
        layer_1_weights[701][4] = 0;
        layer_1_weights[702][4] = 2;
        layer_1_weights[703][4] = -1;
        layer_1_weights[704][4] = 1;
        layer_1_weights[705][4] = 1;
        layer_1_weights[706][4] = 2;
        layer_1_weights[707][4] = 2;
        layer_1_weights[708][4] = 3;
        layer_1_weights[709][4] = 0;
        layer_1_weights[710][4] = 0;
        layer_1_weights[711][4] = -1;
        layer_1_weights[712][4] = -2;
        layer_1_weights[713][4] = 0;
        layer_1_weights[714][4] = 1;
        layer_1_weights[715][4] = 0;
        layer_1_weights[716][4] = -1;
        layer_1_weights[717][4] = 2;
        layer_1_weights[718][4] = 0;
        layer_1_weights[719][4] = 1;
        layer_1_weights[720][4] = -1;
        layer_1_weights[721][4] = -2;
        layer_1_weights[722][4] = -1;
        layer_1_weights[723][4] = 1;
        layer_1_weights[724][4] = -1;
        layer_1_weights[725][4] = 1;
        layer_1_weights[726][4] = -2;
        layer_1_weights[727][4] = 0;
        layer_1_weights[728][4] = 0;
        layer_1_weights[729][4] = 0;
        layer_1_weights[730][4] = 0;
        layer_1_weights[731][4] = 2;
        layer_1_weights[732][4] = 0;
        layer_1_weights[733][4] = 3;
        layer_1_weights[734][4] = 6;
        layer_1_weights[735][4] = 6;
        layer_1_weights[736][4] = 4;
        layer_1_weights[737][4] = 5;
        layer_1_weights[738][4] = 3;
        layer_1_weights[739][4] = -1;
        layer_1_weights[740][4] = 2;
        layer_1_weights[741][4] = 1;
        layer_1_weights[742][4] = 2;
        layer_1_weights[743][4] = 2;
        layer_1_weights[744][4] = 1;
        layer_1_weights[745][4] = 4;
        layer_1_weights[746][4] = 3;
        layer_1_weights[747][4] = 0;
        layer_1_weights[748][4] = 3;
        layer_1_weights[749][4] = 2;
        layer_1_weights[750][4] = -1;
        layer_1_weights[751][4] = 1;
        layer_1_weights[752][4] = 0;
        layer_1_weights[753][4] = -2;
        layer_1_weights[754][4] = 0;
        layer_1_weights[755][4] = 0;
        layer_1_weights[756][4] = 1;
        layer_1_weights[757][4] = 0;
        layer_1_weights[758][4] = 0;
        layer_1_weights[759][4] = 0;
        layer_1_weights[760][4] = -1;
        layer_1_weights[761][4] = -3;
        layer_1_weights[762][4] = 3;
        layer_1_weights[763][4] = 3;
        layer_1_weights[764][4] = 2;
        layer_1_weights[765][4] = 3;
        layer_1_weights[766][4] = 1;
        layer_1_weights[767][4] = 1;
        layer_1_weights[768][4] = 1;
        layer_1_weights[769][4] = 0;
        layer_1_weights[770][4] = 6;
        layer_1_weights[771][4] = 5;
        layer_1_weights[772][4] = 5;
        layer_1_weights[773][4] = 3;
        layer_1_weights[774][4] = 4;
        layer_1_weights[775][4] = 4;
        layer_1_weights[776][4] = 3;
        layer_1_weights[777][4] = 3;
        layer_1_weights[778][4] = 3;
        layer_1_weights[779][4] = 0;
        layer_1_weights[780][4] = 0;
        layer_1_weights[781][4] = 0;
        layer_1_weights[782][4] = 0;
        layer_1_weights[783][4] = 1;
        layer_1_weights[0][5] = 0;
        layer_1_weights[1][5] = 0;
        layer_1_weights[2][5] = 0;
        layer_1_weights[3][5] = 0;
        layer_1_weights[4][5] = 1;
        layer_1_weights[5][5] = -1;
        layer_1_weights[6][5] = 0;
        layer_1_weights[7][5] = 0;
        layer_1_weights[8][5] = 0;
        layer_1_weights[9][5] = 0;
        layer_1_weights[10][5] = 1;
        layer_1_weights[11][5] = 0;
        layer_1_weights[12][5] = 1;
        layer_1_weights[13][5] = 2;
        layer_1_weights[14][5] = 1;
        layer_1_weights[15][5] = 0;
        layer_1_weights[16][5] = 0;
        layer_1_weights[17][5] = 0;
        layer_1_weights[18][5] = -1;
        layer_1_weights[19][5] = 0;
        layer_1_weights[20][5] = 0;
        layer_1_weights[21][5] = 0;
        layer_1_weights[22][5] = -1;
        layer_1_weights[23][5] = 0;
        layer_1_weights[24][5] = 0;
        layer_1_weights[25][5] = 0;
        layer_1_weights[26][5] = 0;
        layer_1_weights[27][5] = 0;
        layer_1_weights[28][5] = 0;
        layer_1_weights[29][5] = 0;
        layer_1_weights[30][5] = 1;
        layer_1_weights[31][5] = 0;
        layer_1_weights[32][5] = 1;
        layer_1_weights[33][5] = 2;
        layer_1_weights[34][5] = -1;
        layer_1_weights[35][5] = -2;
        layer_1_weights[36][5] = -1;
        layer_1_weights[37][5] = -1;
        layer_1_weights[38][5] = -1;
        layer_1_weights[39][5] = -2;
        layer_1_weights[40][5] = -2;
        layer_1_weights[41][5] = 0;
        layer_1_weights[42][5] = -1;
        layer_1_weights[43][5] = 0;
        layer_1_weights[44][5] = -1;
        layer_1_weights[45][5] = -3;
        layer_1_weights[46][5] = 1;
        layer_1_weights[47][5] = 2;
        layer_1_weights[48][5] = 2;
        layer_1_weights[49][5] = -1;
        layer_1_weights[50][5] = 1;
        layer_1_weights[51][5] = 1;
        layer_1_weights[52][5] = 0;
        layer_1_weights[53][5] = 1;
        layer_1_weights[54][5] = 1;
        layer_1_weights[55][5] = 0;
        layer_1_weights[56][5] = 1;
        layer_1_weights[57][5] = 0;
        layer_1_weights[58][5] = 1;
        layer_1_weights[59][5] = 1;
        layer_1_weights[60][5] = 0;
        layer_1_weights[61][5] = -1;
        layer_1_weights[62][5] = -1;
        layer_1_weights[63][5] = 0;
        layer_1_weights[64][5] = 2;
        layer_1_weights[65][5] = 4;
        layer_1_weights[66][5] = 2;
        layer_1_weights[67][5] = 0;
        layer_1_weights[68][5] = 2;
        layer_1_weights[69][5] = 0;
        layer_1_weights[70][5] = 2;
        layer_1_weights[71][5] = 3;
        layer_1_weights[72][5] = 2;
        layer_1_weights[73][5] = 0;
        layer_1_weights[74][5] = 1;
        layer_1_weights[75][5] = -2;
        layer_1_weights[76][5] = 1;
        layer_1_weights[77][5] = 1;
        layer_1_weights[78][5] = -2;
        layer_1_weights[79][5] = 1;
        layer_1_weights[80][5] = 4;
        layer_1_weights[81][5] = 2;
        layer_1_weights[82][5] = 1;
        layer_1_weights[83][5] = 1;
        layer_1_weights[84][5] = 1;
        layer_1_weights[85][5] = 0;
        layer_1_weights[86][5] = 2;
        layer_1_weights[87][5] = 1;
        layer_1_weights[88][5] = -1;
        layer_1_weights[89][5] = 1;
        layer_1_weights[90][5] = 2;
        layer_1_weights[91][5] = 1;
        layer_1_weights[92][5] = 4;
        layer_1_weights[93][5] = 2;
        layer_1_weights[94][5] = 1;
        layer_1_weights[95][5] = -1;
        layer_1_weights[96][5] = 3;
        layer_1_weights[97][5] = 1;
        layer_1_weights[98][5] = 0;
        layer_1_weights[99][5] = 0;
        layer_1_weights[100][5] = 2;
        layer_1_weights[101][5] = 1;
        layer_1_weights[102][5] = 1;
        layer_1_weights[103][5] = 1;
        layer_1_weights[104][5] = 2;
        layer_1_weights[105][5] = 0;
        layer_1_weights[106][5] = 0;
        layer_1_weights[107][5] = -2;
        layer_1_weights[108][5] = -1;
        layer_1_weights[109][5] = -2;
        layer_1_weights[110][5] = -3;
        layer_1_weights[111][5] = 0;
        layer_1_weights[112][5] = 0;
        layer_1_weights[113][5] = 1;
        layer_1_weights[114][5] = 4;
        layer_1_weights[115][5] = 3;
        layer_1_weights[116][5] = 3;
        layer_1_weights[117][5] = 4;
        layer_1_weights[118][5] = 0;
        layer_1_weights[119][5] = -1;
        layer_1_weights[120][5] = 0;
        layer_1_weights[121][5] = -1;
        layer_1_weights[122][5] = -2;
        layer_1_weights[123][5] = -1;
        layer_1_weights[124][5] = -1;
        layer_1_weights[125][5] = 0;
        layer_1_weights[126][5] = -1;
        layer_1_weights[127][5] = 0;
        layer_1_weights[128][5] = 2;
        layer_1_weights[129][5] = 2;
        layer_1_weights[130][5] = -1;
        layer_1_weights[131][5] = 2;
        layer_1_weights[132][5] = 0;
        layer_1_weights[133][5] = 2;
        layer_1_weights[134][5] = 1;
        layer_1_weights[135][5] = -4;
        layer_1_weights[136][5] = -2;
        layer_1_weights[137][5] = -3;
        layer_1_weights[138][5] = 0;
        layer_1_weights[139][5] = -1;
        layer_1_weights[140][5] = 0;
        layer_1_weights[141][5] = 0;
        layer_1_weights[142][5] = 3;
        layer_1_weights[143][5] = -1;
        layer_1_weights[144][5] = 3;
        layer_1_weights[145][5] = 1;
        layer_1_weights[146][5] = 4;
        layer_1_weights[147][5] = 0;
        layer_1_weights[148][5] = -2;
        layer_1_weights[149][5] = 0;
        layer_1_weights[150][5] = -2;
        layer_1_weights[151][5] = -2;
        layer_1_weights[152][5] = -1;
        layer_1_weights[153][5] = -1;
        layer_1_weights[154][5] = 0;
        layer_1_weights[155][5] = 0;
        layer_1_weights[156][5] = 2;
        layer_1_weights[157][5] = 0;
        layer_1_weights[158][5] = 0;
        layer_1_weights[159][5] = -1;
        layer_1_weights[160][5] = 2;
        layer_1_weights[161][5] = 1;
        layer_1_weights[162][5] = 2;
        layer_1_weights[163][5] = 0;
        layer_1_weights[164][5] = 0;
        layer_1_weights[165][5] = 3;
        layer_1_weights[166][5] = 0;
        layer_1_weights[167][5] = -2;
        layer_1_weights[168][5] = 0;
        layer_1_weights[169][5] = 0;
        layer_1_weights[170][5] = 0;
        layer_1_weights[171][5] = 4;
        layer_1_weights[172][5] = 4;
        layer_1_weights[173][5] = 4;
        layer_1_weights[174][5] = 0;
        layer_1_weights[175][5] = 2;
        layer_1_weights[176][5] = 0;
        layer_1_weights[177][5] = 1;
        layer_1_weights[178][5] = 2;
        layer_1_weights[179][5] = 1;
        layer_1_weights[180][5] = 1;
        layer_1_weights[181][5] = -1;
        layer_1_weights[182][5] = -1;
        layer_1_weights[183][5] = -1;
        layer_1_weights[184][5] = 0;
        layer_1_weights[185][5] = -2;
        layer_1_weights[186][5] = -1;
        layer_1_weights[187][5] = 1;
        layer_1_weights[188][5] = 1;
        layer_1_weights[189][5] = 1;
        layer_1_weights[190][5] = 0;
        layer_1_weights[191][5] = 1;
        layer_1_weights[192][5] = 2;
        layer_1_weights[193][5] = 6;
        layer_1_weights[194][5] = 2;
        layer_1_weights[195][5] = 0;
        layer_1_weights[196][5] = -1;
        layer_1_weights[197][5] = 4;
        layer_1_weights[198][5] = 0;
        layer_1_weights[199][5] = 2;
        layer_1_weights[200][5] = 9;
        layer_1_weights[201][5] = 0;
        layer_1_weights[202][5] = 2;
        layer_1_weights[203][5] = 2;
        layer_1_weights[204][5] = -1;
        layer_1_weights[205][5] = 2;
        layer_1_weights[206][5] = 2;
        layer_1_weights[207][5] = 1;
        layer_1_weights[208][5] = 2;
        layer_1_weights[209][5] = 0;
        layer_1_weights[210][5] = -1;
        layer_1_weights[211][5] = 0;
        layer_1_weights[212][5] = -1;
        layer_1_weights[213][5] = 0;
        layer_1_weights[214][5] = 1;
        layer_1_weights[215][5] = 0;
        layer_1_weights[216][5] = 0;
        layer_1_weights[217][5] = 0;
        layer_1_weights[218][5] = 1;
        layer_1_weights[219][5] = 2;
        layer_1_weights[220][5] = -1;
        layer_1_weights[221][5] = 1;
        layer_1_weights[222][5] = -1;
        layer_1_weights[223][5] = 0;
        layer_1_weights[224][5] = 0;
        layer_1_weights[225][5] = 2;
        layer_1_weights[226][5] = 1;
        layer_1_weights[227][5] = 3;
        layer_1_weights[228][5] = 2;
        layer_1_weights[229][5] = 2;
        layer_1_weights[230][5] = 3;
        layer_1_weights[231][5] = 1;
        layer_1_weights[232][5] = 2;
        layer_1_weights[233][5] = 1;
        layer_1_weights[234][5] = 3;
        layer_1_weights[235][5] = 2;
        layer_1_weights[236][5] = 2;
        layer_1_weights[237][5] = 2;
        layer_1_weights[238][5] = 0;
        layer_1_weights[239][5] = 0;
        layer_1_weights[240][5] = 0;
        layer_1_weights[241][5] = 0;
        layer_1_weights[242][5] = -1;
        layer_1_weights[243][5] = 0;
        layer_1_weights[244][5] = 0;
        layer_1_weights[245][5] = -2;
        layer_1_weights[246][5] = 2;
        layer_1_weights[247][5] = -1;
        layer_1_weights[248][5] = 1;
        layer_1_weights[249][5] = 1;
        layer_1_weights[250][5] = 2;
        layer_1_weights[251][5] = 2;
        layer_1_weights[252][5] = 0;
        layer_1_weights[253][5] = 3;
        layer_1_weights[254][5] = 2;
        layer_1_weights[255][5] = 8;
        layer_1_weights[256][5] = 3;
        layer_1_weights[257][5] = 0;
        layer_1_weights[258][5] = 3;
        layer_1_weights[259][5] = 1;
        layer_1_weights[260][5] = 1;
        layer_1_weights[261][5] = 0;
        layer_1_weights[262][5] = 2;
        layer_1_weights[263][5] = 1;
        layer_1_weights[264][5] = 0;
        layer_1_weights[265][5] = 0;
        layer_1_weights[266][5] = 0;
        layer_1_weights[267][5] = 0;
        layer_1_weights[268][5] = 1;
        layer_1_weights[269][5] = 0;
        layer_1_weights[270][5] = 0;
        layer_1_weights[271][5] = 0;
        layer_1_weights[272][5] = 0;
        layer_1_weights[273][5] = 0;
        layer_1_weights[274][5] = 0;
        layer_1_weights[275][5] = 0;
        layer_1_weights[276][5] = 0;
        layer_1_weights[277][5] = -1;
        layer_1_weights[278][5] = 6;
        layer_1_weights[279][5] = 2;
        layer_1_weights[280][5] = 0;
        layer_1_weights[281][5] = 2;
        layer_1_weights[282][5] = 0;
        layer_1_weights[283][5] = 1;
        layer_1_weights[284][5] = 2;
        layer_1_weights[285][5] = -2;
        layer_1_weights[286][5] = 1;
        layer_1_weights[287][5] = 0;
        layer_1_weights[288][5] = 1;
        layer_1_weights[289][5] = -1;
        layer_1_weights[290][5] = 1;
        layer_1_weights[291][5] = -2;
        layer_1_weights[292][5] = -3;
        layer_1_weights[293][5] = -3;
        layer_1_weights[294][5] = 0;
        layer_1_weights[295][5] = -1;
        layer_1_weights[296][5] = -1;
        layer_1_weights[297][5] = 0;
        layer_1_weights[298][5] = 0;
        layer_1_weights[299][5] = 0;
        layer_1_weights[300][5] = 1;
        layer_1_weights[301][5] = -1;
        layer_1_weights[302][5] = 1;
        layer_1_weights[303][5] = -2;
        layer_1_weights[304][5] = -2;
        layer_1_weights[305][5] = 1;
        layer_1_weights[306][5] = 3;
        layer_1_weights[307][5] = 4;
        layer_1_weights[308][5] = 0;
        layer_1_weights[309][5] = 0;
        layer_1_weights[310][5] = -1;
        layer_1_weights[311][5] = 2;
        layer_1_weights[312][5] = 1;
        layer_1_weights[313][5] = -4;
        layer_1_weights[314][5] = -1;
        layer_1_weights[315][5] = 0;
        layer_1_weights[316][5] = -1;
        layer_1_weights[317][5] = -1;
        layer_1_weights[318][5] = -3;
        layer_1_weights[319][5] = -4;
        layer_1_weights[320][5] = -3;
        layer_1_weights[321][5] = -1;
        layer_1_weights[322][5] = 2;
        layer_1_weights[323][5] = 0;
        layer_1_weights[324][5] = -1;
        layer_1_weights[325][5] = -1;
        layer_1_weights[326][5] = -1;
        layer_1_weights[327][5] = -1;
        layer_1_weights[328][5] = 0;
        layer_1_weights[329][5] = -1;
        layer_1_weights[330][5] = -1;
        layer_1_weights[331][5] = 0;
        layer_1_weights[332][5] = -3;
        layer_1_weights[333][5] = 2;
        layer_1_weights[334][5] = 3;
        layer_1_weights[335][5] = 2;
        layer_1_weights[336][5] = 0;
        layer_1_weights[337][5] = -1;
        layer_1_weights[338][5] = 1;
        layer_1_weights[339][5] = -1;
        layer_1_weights[340][5] = -1;
        layer_1_weights[341][5] = -3;
        layer_1_weights[342][5] = -4;
        layer_1_weights[343][5] = -3;
        layer_1_weights[344][5] = -4;
        layer_1_weights[345][5] = -5;
        layer_1_weights[346][5] = -4;
        layer_1_weights[347][5] = -3;
        layer_1_weights[348][5] = -2;
        layer_1_weights[349][5] = 2;
        layer_1_weights[350][5] = 3;
        layer_1_weights[351][5] = 1;
        layer_1_weights[352][5] = 0;
        layer_1_weights[353][5] = 0;
        layer_1_weights[354][5] = -2;
        layer_1_weights[355][5] = 0;
        layer_1_weights[356][5] = -1;
        layer_1_weights[357][5] = 1;
        layer_1_weights[358][5] = -3;
        layer_1_weights[359][5] = -1;
        layer_1_weights[360][5] = -1;
        layer_1_weights[361][5] = 3;
        layer_1_weights[362][5] = 0;
        layer_1_weights[363][5] = 4;
        layer_1_weights[364][5] = 0;
        layer_1_weights[365][5] = -2;
        layer_1_weights[366][5] = -1;
        layer_1_weights[367][5] = 0;
        layer_1_weights[368][5] = -4;
        layer_1_weights[369][5] = -5;
        layer_1_weights[370][5] = -7;
        layer_1_weights[371][5] = -5;
        layer_1_weights[372][5] = -4;
        layer_1_weights[373][5] = -4;
        layer_1_weights[374][5] = -3;
        layer_1_weights[375][5] = -1;
        layer_1_weights[376][5] = 1;
        layer_1_weights[377][5] = 3;
        layer_1_weights[378][5] = 2;
        layer_1_weights[379][5] = 0;
        layer_1_weights[380][5] = 0;
        layer_1_weights[381][5] = -1;
        layer_1_weights[382][5] = -1;
        layer_1_weights[383][5] = 0;
        layer_1_weights[384][5] = 1;
        layer_1_weights[385][5] = 1;
        layer_1_weights[386][5] = -2;
        layer_1_weights[387][5] = 1;
        layer_1_weights[388][5] = 2;
        layer_1_weights[389][5] = 2;
        layer_1_weights[390][5] = 3;
        layer_1_weights[391][5] = 1;
        layer_1_weights[392][5] = -1;
        layer_1_weights[393][5] = 1;
        layer_1_weights[394][5] = 2;
        layer_1_weights[395][5] = -1;
        layer_1_weights[396][5] = -2;
        layer_1_weights[397][5] = -4;
        layer_1_weights[398][5] = -3;
        layer_1_weights[399][5] = -3;
        layer_1_weights[400][5] = -2;
        layer_1_weights[401][5] = -2;
        layer_1_weights[402][5] = 0;
        layer_1_weights[403][5] = 1;
        layer_1_weights[404][5] = 4;
        layer_1_weights[405][5] = 3;
        layer_1_weights[406][5] = 2;
        layer_1_weights[407][5] = 1;
        layer_1_weights[408][5] = -1;
        layer_1_weights[409][5] = -1;
        layer_1_weights[410][5] = 0;
        layer_1_weights[411][5] = 0;
        layer_1_weights[412][5] = -1;
        layer_1_weights[413][5] = 0;
        layer_1_weights[414][5] = 0;
        layer_1_weights[415][5] = 0;
        layer_1_weights[416][5] = 0;
        layer_1_weights[417][5] = 0;
        layer_1_weights[418][5] = 1;
        layer_1_weights[419][5] = -1;
        layer_1_weights[420][5] = 0;
        layer_1_weights[421][5] = 2;
        layer_1_weights[422][5] = 4;
        layer_1_weights[423][5] = 0;
        layer_1_weights[424][5] = -1;
        layer_1_weights[425][5] = 0;
        layer_1_weights[426][5] = 1;
        layer_1_weights[427][5] = -1;
        layer_1_weights[428][5] = -2;
        layer_1_weights[429][5] = 0;
        layer_1_weights[430][5] = 1;
        layer_1_weights[431][5] = 3;
        layer_1_weights[432][5] = 4;
        layer_1_weights[433][5] = 3;
        layer_1_weights[434][5] = 2;
        layer_1_weights[435][5] = 0;
        layer_1_weights[436][5] = -1;
        layer_1_weights[437][5] = -1;
        layer_1_weights[438][5] = 0;
        layer_1_weights[439][5] = 1;
        layer_1_weights[440][5] = -1;
        layer_1_weights[441][5] = 1;
        layer_1_weights[442][5] = 1;
        layer_1_weights[443][5] = -1;
        layer_1_weights[444][5] = 1;
        layer_1_weights[445][5] = -2;
        layer_1_weights[446][5] = 1;
        layer_1_weights[447][5] = 3;
        layer_1_weights[448][5] = 0;
        layer_1_weights[449][5] = 2;
        layer_1_weights[450][5] = 3;
        layer_1_weights[451][5] = 3;
        layer_1_weights[452][5] = 1;
        layer_1_weights[453][5] = 0;
        layer_1_weights[454][5] = 1;
        layer_1_weights[455][5] = 0;
        layer_1_weights[456][5] = 2;
        layer_1_weights[457][5] = 3;
        layer_1_weights[458][5] = 2;
        layer_1_weights[459][5] = 3;
        layer_1_weights[460][5] = 3;
        layer_1_weights[461][5] = 3;
        layer_1_weights[462][5] = 2;
        layer_1_weights[463][5] = 1;
        layer_1_weights[464][5] = 0;
        layer_1_weights[465][5] = 0;
        layer_1_weights[466][5] = 1;
        layer_1_weights[467][5] = 1;
        layer_1_weights[468][5] = 0;
        layer_1_weights[469][5] = 1;
        layer_1_weights[470][5] = 3;
        layer_1_weights[471][5] = 1;
        layer_1_weights[472][5] = 4;
        layer_1_weights[473][5] = -2;
        layer_1_weights[474][5] = 3;
        layer_1_weights[475][5] = 2;
        layer_1_weights[476][5] = 0;
        layer_1_weights[477][5] = 3;
        layer_1_weights[478][5] = 4;
        layer_1_weights[479][5] = 2;
        layer_1_weights[480][5] = 0;
        layer_1_weights[481][5] = 2;
        layer_1_weights[482][5] = 1;
        layer_1_weights[483][5] = 0;
        layer_1_weights[484][5] = 2;
        layer_1_weights[485][5] = 1;
        layer_1_weights[486][5] = 3;
        layer_1_weights[487][5] = 3;
        layer_1_weights[488][5] = 3;
        layer_1_weights[489][5] = 2;
        layer_1_weights[490][5] = 0;
        layer_1_weights[491][5] = 1;
        layer_1_weights[492][5] = 0;
        layer_1_weights[493][5] = 1;
        layer_1_weights[494][5] = 1;
        layer_1_weights[495][5] = 0;
        layer_1_weights[496][5] = 0;
        layer_1_weights[497][5] = -1;
        layer_1_weights[498][5] = 1;
        layer_1_weights[499][5] = 1;
        layer_1_weights[500][5] = 1;
        layer_1_weights[501][5] = -2;
        layer_1_weights[502][5] = 3;
        layer_1_weights[503][5] = -2;
        layer_1_weights[504][5] = -1;
        layer_1_weights[505][5] = 0;
        layer_1_weights[506][5] = 3;
        layer_1_weights[507][5] = 5;
        layer_1_weights[508][5] = 1;
        layer_1_weights[509][5] = 2;
        layer_1_weights[510][5] = 0;
        layer_1_weights[511][5] = 0;
        layer_1_weights[512][5] = 2;
        layer_1_weights[513][5] = 2;
        layer_1_weights[514][5] = 2;
        layer_1_weights[515][5] = 1;
        layer_1_weights[516][5] = 1;
        layer_1_weights[517][5] = 0;
        layer_1_weights[518][5] = 0;
        layer_1_weights[519][5] = 0;
        layer_1_weights[520][5] = 1;
        layer_1_weights[521][5] = 0;
        layer_1_weights[522][5] = 1;
        layer_1_weights[523][5] = 0;
        layer_1_weights[524][5] = -1;
        layer_1_weights[525][5] = 1;
        layer_1_weights[526][5] = -1;
        layer_1_weights[527][5] = 2;
        layer_1_weights[528][5] = 1;
        layer_1_weights[529][5] = 1;
        layer_1_weights[530][5] = 5;
        layer_1_weights[531][5] = 3;
        layer_1_weights[532][5] = 1;
        layer_1_weights[533][5] = -2;
        layer_1_weights[534][5] = 0;
        layer_1_weights[535][5] = 2;
        layer_1_weights[536][5] = 3;
        layer_1_weights[537][5] = 1;
        layer_1_weights[538][5] = 1;
        layer_1_weights[539][5] = 1;
        layer_1_weights[540][5] = 2;
        layer_1_weights[541][5] = 3;
        layer_1_weights[542][5] = 1;
        layer_1_weights[543][5] = 1;
        layer_1_weights[544][5] = 1;
        layer_1_weights[545][5] = -1;
        layer_1_weights[546][5] = -1;
        layer_1_weights[547][5] = 0;
        layer_1_weights[548][5] = -1;
        layer_1_weights[549][5] = 0;
        layer_1_weights[550][5] = 0;
        layer_1_weights[551][5] = 0;
        layer_1_weights[552][5] = -1;
        layer_1_weights[553][5] = 0;
        layer_1_weights[554][5] = 1;
        layer_1_weights[555][5] = 1;
        layer_1_weights[556][5] = -2;
        layer_1_weights[557][5] = 0;
        layer_1_weights[558][5] = 3;
        layer_1_weights[559][5] = 3;
        layer_1_weights[560][5] = 0;
        layer_1_weights[561][5] = -1;
        layer_1_weights[562][5] = 0;
        layer_1_weights[563][5] = 2;
        layer_1_weights[564][5] = -1;
        layer_1_weights[565][5] = -2;
        layer_1_weights[566][5] = 2;
        layer_1_weights[567][5] = 3;
        layer_1_weights[568][5] = 0;
        layer_1_weights[569][5] = 1;
        layer_1_weights[570][5] = 0;
        layer_1_weights[571][5] = -1;
        layer_1_weights[572][5] = 1;
        layer_1_weights[573][5] = -1;
        layer_1_weights[574][5] = -1;
        layer_1_weights[575][5] = -1;
        layer_1_weights[576][5] = -1;
        layer_1_weights[577][5] = -1;
        layer_1_weights[578][5] = -1;
        layer_1_weights[579][5] = -1;
        layer_1_weights[580][5] = 0;
        layer_1_weights[581][5] = 1;
        layer_1_weights[582][5] = 0;
        layer_1_weights[583][5] = 1;
        layer_1_weights[584][5] = -2;
        layer_1_weights[585][5] = -2;
        layer_1_weights[586][5] = 2;
        layer_1_weights[587][5] = 1;
        layer_1_weights[588][5] = 1;
        layer_1_weights[589][5] = 3;
        layer_1_weights[590][5] = 6;
        layer_1_weights[591][5] = -1;
        layer_1_weights[592][5] = 1;
        layer_1_weights[593][5] = 0;
        layer_1_weights[594][5] = 4;
        layer_1_weights[595][5] = 1;
        layer_1_weights[596][5] = -1;
        layer_1_weights[597][5] = 2;
        layer_1_weights[598][5] = 0;
        layer_1_weights[599][5] = 0;
        layer_1_weights[600][5] = 1;
        layer_1_weights[601][5] = 0;
        layer_1_weights[602][5] = 0;
        layer_1_weights[603][5] = -1;
        layer_1_weights[604][5] = 0;
        layer_1_weights[605][5] = -1;
        layer_1_weights[606][5] = -1;
        layer_1_weights[607][5] = -2;
        layer_1_weights[608][5] = 1;
        layer_1_weights[609][5] = -1;
        layer_1_weights[610][5] = 1;
        layer_1_weights[611][5] = 0;
        layer_1_weights[612][5] = -4;
        layer_1_weights[613][5] = -4;
        layer_1_weights[614][5] = -2;
        layer_1_weights[615][5] = 0;
        layer_1_weights[616][5] = 0;
        layer_1_weights[617][5] = 2;
        layer_1_weights[618][5] = 3;
        layer_1_weights[619][5] = 2;
        layer_1_weights[620][5] = 3;
        layer_1_weights[621][5] = 1;
        layer_1_weights[622][5] = 0;
        layer_1_weights[623][5] = 2;
        layer_1_weights[624][5] = -1;
        layer_1_weights[625][5] = 0;
        layer_1_weights[626][5] = 1;
        layer_1_weights[627][5] = 0;
        layer_1_weights[628][5] = -1;
        layer_1_weights[629][5] = -1;
        layer_1_weights[630][5] = 0;
        layer_1_weights[631][5] = 0;
        layer_1_weights[632][5] = -1;
        layer_1_weights[633][5] = 0;
        layer_1_weights[634][5] = -2;
        layer_1_weights[635][5] = 0;
        layer_1_weights[636][5] = 0;
        layer_1_weights[637][5] = -1;
        layer_1_weights[638][5] = -1;
        layer_1_weights[639][5] = -1;
        layer_1_weights[640][5] = -4;
        layer_1_weights[641][5] = -3;
        layer_1_weights[642][5] = -3;
        layer_1_weights[643][5] = 0;
        layer_1_weights[644][5] = 0;
        layer_1_weights[645][5] = 0;
        layer_1_weights[646][5] = 2;
        layer_1_weights[647][5] = -1;
        layer_1_weights[648][5] = 4;
        layer_1_weights[649][5] = 0;
        layer_1_weights[650][5] = 2;
        layer_1_weights[651][5] = 0;
        layer_1_weights[652][5] = -1;
        layer_1_weights[653][5] = 0;
        layer_1_weights[654][5] = -2;
        layer_1_weights[655][5] = 0;
        layer_1_weights[656][5] = 0;
        layer_1_weights[657][5] = 1;
        layer_1_weights[658][5] = 1;
        layer_1_weights[659][5] = 0;
        layer_1_weights[660][5] = 0;
        layer_1_weights[661][5] = 0;
        layer_1_weights[662][5] = 0;
        layer_1_weights[663][5] = 0;
        layer_1_weights[664][5] = -2;
        layer_1_weights[665][5] = 0;
        layer_1_weights[666][5] = -1;
        layer_1_weights[667][5] = -2;
        layer_1_weights[668][5] = -5;
        layer_1_weights[669][5] = -4;
        layer_1_weights[670][5] = -1;
        layer_1_weights[671][5] = 0;
        layer_1_weights[672][5] = 0;
        layer_1_weights[673][5] = 0;
        layer_1_weights[674][5] = 3;
        layer_1_weights[675][5] = 0;
        layer_1_weights[676][5] = 1;
        layer_1_weights[677][5] = 0;
        layer_1_weights[678][5] = 1;
        layer_1_weights[679][5] = 0;
        layer_1_weights[680][5] = 0;
        layer_1_weights[681][5] = 2;
        layer_1_weights[682][5] = 0;
        layer_1_weights[683][5] = 1;
        layer_1_weights[684][5] = 0;
        layer_1_weights[685][5] = 0;
        layer_1_weights[686][5] = 0;
        layer_1_weights[687][5] = -1;
        layer_1_weights[688][5] = -1;
        layer_1_weights[689][5] = 0;
        layer_1_weights[690][5] = -4;
        layer_1_weights[691][5] = -2;
        layer_1_weights[692][5] = -1;
        layer_1_weights[693][5] = -4;
        layer_1_weights[694][5] = -4;
        layer_1_weights[695][5] = -5;
        layer_1_weights[696][5] = -4;
        layer_1_weights[697][5] = 0;
        layer_1_weights[698][5] = 2;
        layer_1_weights[699][5] = 0;
        layer_1_weights[700][5] = 0;
        layer_1_weights[701][5] = 0;
        layer_1_weights[702][5] = -1;
        layer_1_weights[703][5] = 0;
        layer_1_weights[704][5] = -2;
        layer_1_weights[705][5] = 0;
        layer_1_weights[706][5] = 1;
        layer_1_weights[707][5] = 0;
        layer_1_weights[708][5] = -1;
        layer_1_weights[709][5] = 1;
        layer_1_weights[710][5] = 0;
        layer_1_weights[711][5] = 1;
        layer_1_weights[712][5] = 1;
        layer_1_weights[713][5] = 1;
        layer_1_weights[714][5] = 0;
        layer_1_weights[715][5] = -1;
        layer_1_weights[716][5] = 0;
        layer_1_weights[717][5] = -1;
        layer_1_weights[718][5] = -1;
        layer_1_weights[719][5] = 0;
        layer_1_weights[720][5] = 0;
        layer_1_weights[721][5] = -2;
        layer_1_weights[722][5] = -5;
        layer_1_weights[723][5] = -4;
        layer_1_weights[724][5] = -4;
        layer_1_weights[725][5] = -1;
        layer_1_weights[726][5] = 2;
        layer_1_weights[727][5] = 1;
        layer_1_weights[728][5] = 0;
        layer_1_weights[729][5] = 0;
        layer_1_weights[730][5] = -1;
        layer_1_weights[731][5] = -2;
        layer_1_weights[732][5] = -2;
        layer_1_weights[733][5] = 0;
        layer_1_weights[734][5] = -2;
        layer_1_weights[735][5] = 0;
        layer_1_weights[736][5] = 0;
        layer_1_weights[737][5] = -1;
        layer_1_weights[738][5] = 1;
        layer_1_weights[739][5] = -1;
        layer_1_weights[740][5] = -3;
        layer_1_weights[741][5] = -1;
        layer_1_weights[742][5] = -3;
        layer_1_weights[743][5] = -3;
        layer_1_weights[744][5] = -2;
        layer_1_weights[745][5] = -4;
        layer_1_weights[746][5] = -2;
        layer_1_weights[747][5] = -1;
        layer_1_weights[748][5] = -1;
        layer_1_weights[749][5] = -4;
        layer_1_weights[750][5] = -3;
        layer_1_weights[751][5] = 0;
        layer_1_weights[752][5] = 0;
        layer_1_weights[753][5] = 3;
        layer_1_weights[754][5] = 0;
        layer_1_weights[755][5] = 0;
        layer_1_weights[756][5] = 0;
        layer_1_weights[757][5] = 0;
        layer_1_weights[758][5] = 0;
        layer_1_weights[759][5] = 1;
        layer_1_weights[760][5] = 1;
        layer_1_weights[761][5] = 2;
        layer_1_weights[762][5] = 2;
        layer_1_weights[763][5] = 3;
        layer_1_weights[764][5] = 1;
        layer_1_weights[765][5] = 2;
        layer_1_weights[766][5] = 6;
        layer_1_weights[767][5] = 3;
        layer_1_weights[768][5] = -1;
        layer_1_weights[769][5] = -2;
        layer_1_weights[770][5] = -1;
        layer_1_weights[771][5] = 0;
        layer_1_weights[772][5] = 3;
        layer_1_weights[773][5] = 1;
        layer_1_weights[774][5] = 0;
        layer_1_weights[775][5] = 2;
        layer_1_weights[776][5] = -1;
        layer_1_weights[777][5] = 0;
        layer_1_weights[778][5] = -2;
        layer_1_weights[779][5] = 1;
        layer_1_weights[780][5] = -1;
        layer_1_weights[781][5] = 0;
        layer_1_weights[782][5] = 0;
        layer_1_weights[783][5] = 1;
        layer_1_weights[0][6] = 0;
        layer_1_weights[1][6] = 0;
        layer_1_weights[2][6] = 0;
        layer_1_weights[3][6] = -1;
        layer_1_weights[4][6] = 0;
        layer_1_weights[5][6] = 0;
        layer_1_weights[6][6] = 0;
        layer_1_weights[7][6] = -1;
        layer_1_weights[8][6] = 0;
        layer_1_weights[9][6] = 1;
        layer_1_weights[10][6] = -1;
        layer_1_weights[11][6] = 0;
        layer_1_weights[12][6] = -1;
        layer_1_weights[13][6] = 2;
        layer_1_weights[14][6] = 2;
        layer_1_weights[15][6] = 0;
        layer_1_weights[16][6] = 0;
        layer_1_weights[17][6] = 0;
        layer_1_weights[18][6] = 0;
        layer_1_weights[19][6] = -1;
        layer_1_weights[20][6] = 0;
        layer_1_weights[21][6] = 0;
        layer_1_weights[22][6] = 0;
        layer_1_weights[23][6] = 0;
        layer_1_weights[24][6] = 0;
        layer_1_weights[25][6] = 0;
        layer_1_weights[26][6] = 1;
        layer_1_weights[27][6] = 0;
        layer_1_weights[28][6] = 0;
        layer_1_weights[29][6] = 0;
        layer_1_weights[30][6] = 0;
        layer_1_weights[31][6] = 0;
        layer_1_weights[32][6] = 0;
        layer_1_weights[33][6] = -1;
        layer_1_weights[34][6] = 0;
        layer_1_weights[35][6] = -2;
        layer_1_weights[36][6] = 0;
        layer_1_weights[37][6] = -1;
        layer_1_weights[38][6] = -1;
        layer_1_weights[39][6] = 1;
        layer_1_weights[40][6] = -3;
        layer_1_weights[41][6] = -2;
        layer_1_weights[42][6] = -2;
        layer_1_weights[43][6] = 1;
        layer_1_weights[44][6] = 1;
        layer_1_weights[45][6] = 0;
        layer_1_weights[46][6] = -1;
        layer_1_weights[47][6] = -5;
        layer_1_weights[48][6] = -5;
        layer_1_weights[49][6] = -4;
        layer_1_weights[50][6] = -2;
        layer_1_weights[51][6] = 0;
        layer_1_weights[52][6] = 0;
        layer_1_weights[53][6] = 1;
        layer_1_weights[54][6] = 0;
        layer_1_weights[55][6] = 1;
        layer_1_weights[56][6] = 0;
        layer_1_weights[57][6] = 0;
        layer_1_weights[58][6] = -1;
        layer_1_weights[59][6] = 0;
        layer_1_weights[60][6] = -2;
        layer_1_weights[61][6] = 1;
        layer_1_weights[62][6] = 1;
        layer_1_weights[63][6] = 1;
        layer_1_weights[64][6] = 2;
        layer_1_weights[65][6] = 3;
        layer_1_weights[66][6] = 0;
        layer_1_weights[67][6] = -2;
        layer_1_weights[68][6] = 1;
        layer_1_weights[69][6] = -2;
        layer_1_weights[70][6] = 1;
        layer_1_weights[71][6] = 0;
        layer_1_weights[72][6] = 3;
        layer_1_weights[73][6] = 0;
        layer_1_weights[74][6] = 1;
        layer_1_weights[75][6] = 0;
        layer_1_weights[76][6] = 0;
        layer_1_weights[77][6] = 0;
        layer_1_weights[78][6] = -1;
        layer_1_weights[79][6] = 1;
        layer_1_weights[80][6] = 0;
        layer_1_weights[81][6] = -1;
        layer_1_weights[82][6] = 0;
        layer_1_weights[83][6] = 0;
        layer_1_weights[84][6] = 0;
        layer_1_weights[85][6] = 0;
        layer_1_weights[86][6] = 2;
        layer_1_weights[87][6] = 0;
        layer_1_weights[88][6] = 3;
        layer_1_weights[89][6] = -2;
        layer_1_weights[90][6] = 1;
        layer_1_weights[91][6] = 1;
        layer_1_weights[92][6] = 2;
        layer_1_weights[93][6] = 2;
        layer_1_weights[94][6] = 1;
        layer_1_weights[95][6] = -1;
        layer_1_weights[96][6] = -1;
        layer_1_weights[97][6] = -1;
        layer_1_weights[98][6] = -2;
        layer_1_weights[99][6] = -1;
        layer_1_weights[100][6] = 0;
        layer_1_weights[101][6] = 0;
        layer_1_weights[102][6] = 0;
        layer_1_weights[103][6] = 2;
        layer_1_weights[104][6] = 0;
        layer_1_weights[105][6] = 0;
        layer_1_weights[106][6] = 0;
        layer_1_weights[107][6] = -4;
        layer_1_weights[108][6] = 1;
        layer_1_weights[109][6] = -1;
        layer_1_weights[110][6] = 0;
        layer_1_weights[111][6] = 0;
        layer_1_weights[112][6] = 0;
        layer_1_weights[113][6] = -2;
        layer_1_weights[114][6] = 1;
        layer_1_weights[115][6] = -3;
        layer_1_weights[116][6] = 0;
        layer_1_weights[117][6] = 0;
        layer_1_weights[118][6] = 0;
        layer_1_weights[119][6] = 2;
        layer_1_weights[120][6] = 0;
        layer_1_weights[121][6] = 1;
        layer_1_weights[122][6] = 0;
        layer_1_weights[123][6] = 1;
        layer_1_weights[124][6] = 1;
        layer_1_weights[125][6] = 0;
        layer_1_weights[126][6] = -1;
        layer_1_weights[127][6] = -1;
        layer_1_weights[128][6] = 0;
        layer_1_weights[129][6] = 0;
        layer_1_weights[130][6] = 1;
        layer_1_weights[131][6] = -1;
        layer_1_weights[132][6] = -2;
        layer_1_weights[133][6] = -2;
        layer_1_weights[134][6] = -2;
        layer_1_weights[135][6] = 0;
        layer_1_weights[136][6] = -1;
        layer_1_weights[137][6] = -2;
        layer_1_weights[138][6] = -2;
        layer_1_weights[139][6] = -2;
        layer_1_weights[140][6] = 0;
        layer_1_weights[141][6] = 0;
        layer_1_weights[142][6] = 0;
        layer_1_weights[143][6] = 3;
        layer_1_weights[144][6] = 2;
        layer_1_weights[145][6] = 0;
        layer_1_weights[146][6] = 0;
        layer_1_weights[147][6] = -3;
        layer_1_weights[148][6] = -3;
        layer_1_weights[149][6] = -1;
        layer_1_weights[150][6] = 0;
        layer_1_weights[151][6] = 2;
        layer_1_weights[152][6] = 0;
        layer_1_weights[153][6] = 0;
        layer_1_weights[154][6] = -1;
        layer_1_weights[155][6] = 0;
        layer_1_weights[156][6] = -1;
        layer_1_weights[157][6] = -1;
        layer_1_weights[158][6] = 0;
        layer_1_weights[159][6] = -1;
        layer_1_weights[160][6] = 0;
        layer_1_weights[161][6] = 1;
        layer_1_weights[162][6] = 2;
        layer_1_weights[163][6] = 0;
        layer_1_weights[164][6] = -1;
        layer_1_weights[165][6] = 0;
        layer_1_weights[166][6] = 0;
        layer_1_weights[167][6] = -2;
        layer_1_weights[168][6] = 0;
        layer_1_weights[169][6] = 0;
        layer_1_weights[170][6] = 1;
        layer_1_weights[171][6] = -1;
        layer_1_weights[172][6] = 0;
        layer_1_weights[173][6] = -3;
        layer_1_weights[174][6] = -1;
        layer_1_weights[175][6] = -3;
        layer_1_weights[176][6] = 0;
        layer_1_weights[177][6] = -2;
        layer_1_weights[178][6] = 1;
        layer_1_weights[179][6] = 1;
        layer_1_weights[180][6] = 0;
        layer_1_weights[181][6] = 0;
        layer_1_weights[182][6] = 1;
        layer_1_weights[183][6] = -1;
        layer_1_weights[184][6] = 0;
        layer_1_weights[185][6] = -1;
        layer_1_weights[186][6] = 0;
        layer_1_weights[187][6] = 0;
        layer_1_weights[188][6] = 1;
        layer_1_weights[189][6] = 0;
        layer_1_weights[190][6] = 0;
        layer_1_weights[191][6] = 1;
        layer_1_weights[192][6] = 1;
        layer_1_weights[193][6] = 0;
        layer_1_weights[194][6] = 1;
        layer_1_weights[195][6] = -1;
        layer_1_weights[196][6] = -1;
        layer_1_weights[197][6] = -2;
        layer_1_weights[198][6] = 1;
        layer_1_weights[199][6] = -1;
        layer_1_weights[200][6] = -5;
        layer_1_weights[201][6] = -4;
        layer_1_weights[202][6] = -1;
        layer_1_weights[203][6] = -1;
        layer_1_weights[204][6] = 0;
        layer_1_weights[205][6] = -1;
        layer_1_weights[206][6] = 0;
        layer_1_weights[207][6] = 1;
        layer_1_weights[208][6] = 1;
        layer_1_weights[209][6] = 2;
        layer_1_weights[210][6] = 1;
        layer_1_weights[211][6] = 0;
        layer_1_weights[212][6] = 0;
        layer_1_weights[213][6] = -1;
        layer_1_weights[214][6] = 0;
        layer_1_weights[215][6] = -1;
        layer_1_weights[216][6] = -1;
        layer_1_weights[217][6] = 0;
        layer_1_weights[218][6] = 2;
        layer_1_weights[219][6] = 0;
        layer_1_weights[220][6] = 1;
        layer_1_weights[221][6] = 0;
        layer_1_weights[222][6] = 0;
        layer_1_weights[223][6] = 0;
        layer_1_weights[224][6] = 0;
        layer_1_weights[225][6] = 2;
        layer_1_weights[226][6] = -1;
        layer_1_weights[227][6] = -4;
        layer_1_weights[228][6] = -5;
        layer_1_weights[229][6] = 0;
        layer_1_weights[230][6] = -3;
        layer_1_weights[231][6] = -1;
        layer_1_weights[232][6] = -2;
        layer_1_weights[233][6] = -1;
        layer_1_weights[234][6] = -1;
        layer_1_weights[235][6] = 0;
        layer_1_weights[236][6] = 2;
        layer_1_weights[237][6] = 1;
        layer_1_weights[238][6] = 2;
        layer_1_weights[239][6] = 1;
        layer_1_weights[240][6] = 0;
        layer_1_weights[241][6] = 1;
        layer_1_weights[242][6] = 1;
        layer_1_weights[243][6] = 1;
        layer_1_weights[244][6] = 0;
        layer_1_weights[245][6] = 0;
        layer_1_weights[246][6] = 0;
        layer_1_weights[247][6] = 1;
        layer_1_weights[248][6] = 1;
        layer_1_weights[249][6] = 0;
        layer_1_weights[250][6] = -1;
        layer_1_weights[251][6] = 3;
        layer_1_weights[252][6] = -2;
        layer_1_weights[253][6] = -2;
        layer_1_weights[254][6] = -5;
        layer_1_weights[255][6] = 1;
        layer_1_weights[256][6] = -4;
        layer_1_weights[257][6] = -1;
        layer_1_weights[258][6] = -3;
        layer_1_weights[259][6] = -2;
        layer_1_weights[260][6] = -1;
        layer_1_weights[261][6] = 0;
        layer_1_weights[262][6] = 0;
        layer_1_weights[263][6] = 0;
        layer_1_weights[264][6] = 1;
        layer_1_weights[265][6] = 1;
        layer_1_weights[266][6] = 2;
        layer_1_weights[267][6] = 3;
        layer_1_weights[268][6] = 1;
        layer_1_weights[269][6] = 1;
        layer_1_weights[270][6] = 1;
        layer_1_weights[271][6] = 0;
        layer_1_weights[272][6] = -1;
        layer_1_weights[273][6] = -1;
        layer_1_weights[274][6] = 1;
        layer_1_weights[275][6] = 2;
        layer_1_weights[276][6] = 0;
        layer_1_weights[277][6] = 3;
        layer_1_weights[278][6] = 1;
        layer_1_weights[279][6] = -2;
        layer_1_weights[280][6] = -2;
        layer_1_weights[281][6] = 0;
        layer_1_weights[282][6] = 0;
        layer_1_weights[283][6] = 1;
        layer_1_weights[284][6] = -2;
        layer_1_weights[285][6] = 0;
        layer_1_weights[286][6] = 1;
        layer_1_weights[287][6] = 1;
        layer_1_weights[288][6] = 1;
        layer_1_weights[289][6] = 0;
        layer_1_weights[290][6] = 1;
        layer_1_weights[291][6] = 1;
        layer_1_weights[292][6] = 0;
        layer_1_weights[293][6] = 1;
        layer_1_weights[294][6] = 1;
        layer_1_weights[295][6] = 2;
        layer_1_weights[296][6] = 1;
        layer_1_weights[297][6] = 0;
        layer_1_weights[298][6] = 0;
        layer_1_weights[299][6] = 0;
        layer_1_weights[300][6] = -2;
        layer_1_weights[301][6] = 1;
        layer_1_weights[302][6] = -1;
        layer_1_weights[303][6] = 2;
        layer_1_weights[304][6] = 1;
        layer_1_weights[305][6] = 4;
        layer_1_weights[306][6] = 5;
        layer_1_weights[307][6] = 0;
        layer_1_weights[308][6] = -3;
        layer_1_weights[309][6] = 2;
        layer_1_weights[310][6] = 0;
        layer_1_weights[311][6] = -1;
        layer_1_weights[312][6] = 1;
        layer_1_weights[313][6] = 3;
        layer_1_weights[314][6] = 0;
        layer_1_weights[315][6] = -1;
        layer_1_weights[316][6] = -2;
        layer_1_weights[317][6] = -2;
        layer_1_weights[318][6] = -1;
        layer_1_weights[319][6] = 0;
        layer_1_weights[320][6] = -1;
        layer_1_weights[321][6] = -2;
        layer_1_weights[322][6] = 0;
        layer_1_weights[323][6] = 1;
        layer_1_weights[324][6] = 0;
        layer_1_weights[325][6] = 0;
        layer_1_weights[326][6] = 0;
        layer_1_weights[327][6] = 1;
        layer_1_weights[328][6] = 0;
        layer_1_weights[329][6] = -1;
        layer_1_weights[330][6] = 2;
        layer_1_weights[331][6] = -1;
        layer_1_weights[332][6] = 3;
        layer_1_weights[333][6] = 6;
        layer_1_weights[334][6] = 1;
        layer_1_weights[335][6] = 1;
        layer_1_weights[336][6] = -2;
        layer_1_weights[337][6] = -3;
        layer_1_weights[338][6] = -2;
        layer_1_weights[339][6] = 2;
        layer_1_weights[340][6] = 0;
        layer_1_weights[341][6] = 1;
        layer_1_weights[342][6] = -1;
        layer_1_weights[343][6] = 0;
        layer_1_weights[344][6] = -1;
        layer_1_weights[345][6] = -1;
        layer_1_weights[346][6] = -2;
        layer_1_weights[347][6] = -2;
        layer_1_weights[348][6] = -2;
        layer_1_weights[349][6] = 0;
        layer_1_weights[350][6] = 1;
        layer_1_weights[351][6] = 0;
        layer_1_weights[352][6] = -1;
        layer_1_weights[353][6] = -1;
        layer_1_weights[354][6] = 0;
        layer_1_weights[355][6] = 0;
        layer_1_weights[356][6] = -1;
        layer_1_weights[357][6] = -1;
        layer_1_weights[358][6] = -2;
        layer_1_weights[359][6] = -3;
        layer_1_weights[360][6] = -4;
        layer_1_weights[361][6] = 0;
        layer_1_weights[362][6] = 3;
        layer_1_weights[363][6] = -1;
        layer_1_weights[364][6] = 0;
        layer_1_weights[365][6] = -1;
        layer_1_weights[366][6] = -1;
        layer_1_weights[367][6] = 3;
        layer_1_weights[368][6] = 0;
        layer_1_weights[369][6] = 0;
        layer_1_weights[370][6] = -1;
        layer_1_weights[371][6] = 0;
        layer_1_weights[372][6] = 0;
        layer_1_weights[373][6] = -1;
        layer_1_weights[374][6] = -2;
        layer_1_weights[375][6] = -1;
        layer_1_weights[376][6] = 2;
        layer_1_weights[377][6] = 3;
        layer_1_weights[378][6] = 2;
        layer_1_weights[379][6] = 0;
        layer_1_weights[380][6] = -2;
        layer_1_weights[381][6] = 0;
        layer_1_weights[382][6] = -2;
        layer_1_weights[383][6] = -1;
        layer_1_weights[384][6] = -1;
        layer_1_weights[385][6] = -1;
        layer_1_weights[386][6] = -1;
        layer_1_weights[387][6] = -1;
        layer_1_weights[388][6] = -2;
        layer_1_weights[389][6] = -1;
        layer_1_weights[390][6] = 5;
        layer_1_weights[391][6] = 0;
        layer_1_weights[392][6] = 3;
        layer_1_weights[393][6] = -2;
        layer_1_weights[394][6] = -3;
        layer_1_weights[395][6] = 2;
        layer_1_weights[396][6] = -2;
        layer_1_weights[397][6] = -2;
        layer_1_weights[398][6] = 0;
        layer_1_weights[399][6] = 0;
        layer_1_weights[400][6] = -2;
        layer_1_weights[401][6] = -1;
        layer_1_weights[402][6] = 0;
        layer_1_weights[403][6] = -1;
        layer_1_weights[404][6] = 1;
        layer_1_weights[405][6] = 3;
        layer_1_weights[406][6] = 0;
        layer_1_weights[407][6] = 0;
        layer_1_weights[408][6] = 0;
        layer_1_weights[409][6] = 0;
        layer_1_weights[410][6] = 0;
        layer_1_weights[411][6] = -1;
        layer_1_weights[412][6] = 0;
        layer_1_weights[413][6] = -1;
        layer_1_weights[414][6] = -2;
        layer_1_weights[415][6] = -2;
        layer_1_weights[416][6] = 0;
        layer_1_weights[417][6] = -2;
        layer_1_weights[418][6] = 2;
        layer_1_weights[419][6] = 2;
        layer_1_weights[420][6] = 2;
        layer_1_weights[421][6] = -2;
        layer_1_weights[422][6] = -3;
        layer_1_weights[423][6] = 1;
        layer_1_weights[424][6] = 1;
        layer_1_weights[425][6] = 1;
        layer_1_weights[426][6] = 0;
        layer_1_weights[427][6] = -1;
        layer_1_weights[428][6] = -1;
        layer_1_weights[429][6] = 0;
        layer_1_weights[430][6] = 0;
        layer_1_weights[431][6] = 1;
        layer_1_weights[432][6] = 2;
        layer_1_weights[433][6] = 2;
        layer_1_weights[434][6] = 1;
        layer_1_weights[435][6] = -1;
        layer_1_weights[436][6] = 0;
        layer_1_weights[437][6] = -1;
        layer_1_weights[438][6] = 0;
        layer_1_weights[439][6] = -1;
        layer_1_weights[440][6] = -2;
        layer_1_weights[441][6] = -2;
        layer_1_weights[442][6] = -3;
        layer_1_weights[443][6] = -3;
        layer_1_weights[444][6] = 1;
        layer_1_weights[445][6] = 1;
        layer_1_weights[446][6] = 4;
        layer_1_weights[447][6] = 3;
        layer_1_weights[448][6] = -2;
        layer_1_weights[449][6] = -1;
        layer_1_weights[450][6] = 1;
        layer_1_weights[451][6] = 2;
        layer_1_weights[452][6] = 0;
        layer_1_weights[453][6] = 1;
        layer_1_weights[454][6] = 1;
        layer_1_weights[455][6] = -1;
        layer_1_weights[456][6] = -1;
        layer_1_weights[457][6] = 0;
        layer_1_weights[458][6] = 0;
        layer_1_weights[459][6] = 0;
        layer_1_weights[460][6] = 1;
        layer_1_weights[461][6] = 1;
        layer_1_weights[462][6] = 1;
        layer_1_weights[463][6] = 0;
        layer_1_weights[464][6] = 1;
        layer_1_weights[465][6] = 0;
        layer_1_weights[466][6] = -1;
        layer_1_weights[467][6] = -3;
        layer_1_weights[468][6] = -1;
        layer_1_weights[469][6] = -1;
        layer_1_weights[470][6] = 0;
        layer_1_weights[471][6] = -1;
        layer_1_weights[472][6] = -1;
        layer_1_weights[473][6] = 2;
        layer_1_weights[474][6] = 3;
        layer_1_weights[475][6] = 4;
        layer_1_weights[476][6] = 0;
        layer_1_weights[477][6] = -1;
        layer_1_weights[478][6] = -2;
        layer_1_weights[479][6] = 2;
        layer_1_weights[480][6] = 1;
        layer_1_weights[481][6] = 2;
        layer_1_weights[482][6] = 2;
        layer_1_weights[483][6] = 1;
        layer_1_weights[484][6] = 0;
        layer_1_weights[485][6] = 1;
        layer_1_weights[486][6] = 1;
        layer_1_weights[487][6] = 1;
        layer_1_weights[488][6] = 0;
        layer_1_weights[489][6] = 1;
        layer_1_weights[490][6] = 2;
        layer_1_weights[491][6] = 0;
        layer_1_weights[492][6] = 0;
        layer_1_weights[493][6] = 0;
        layer_1_weights[494][6] = 0;
        layer_1_weights[495][6] = -1;
        layer_1_weights[496][6] = -1;
        layer_1_weights[497][6] = -1;
        layer_1_weights[498][6] = -1;
        layer_1_weights[499][6] = -1;
        layer_1_weights[500][6] = -1;
        layer_1_weights[501][6] = 2;
        layer_1_weights[502][6] = 1;
        layer_1_weights[503][6] = 5;
        layer_1_weights[504][6] = 2;
        layer_1_weights[505][6] = -1;
        layer_1_weights[506][6] = -2;
        layer_1_weights[507][6] = -1;
        layer_1_weights[508][6] = 3;
        layer_1_weights[509][6] = 2;
        layer_1_weights[510][6] = 2;
        layer_1_weights[511][6] = 1;
        layer_1_weights[512][6] = 0;
        layer_1_weights[513][6] = 1;
        layer_1_weights[514][6] = 0;
        layer_1_weights[515][6] = 0;
        layer_1_weights[516][6] = 1;
        layer_1_weights[517][6] = 1;
        layer_1_weights[518][6] = 1;
        layer_1_weights[519][6] = 1;
        layer_1_weights[520][6] = 1;
        layer_1_weights[521][6] = 1;
        layer_1_weights[522][6] = -1;
        layer_1_weights[523][6] = -1;
        layer_1_weights[524][6] = 0;
        layer_1_weights[525][6] = -1;
        layer_1_weights[526][6] = 0;
        layer_1_weights[527][6] = 0;
        layer_1_weights[528][6] = 2;
        layer_1_weights[529][6] = 4;
        layer_1_weights[530][6] = -1;
        layer_1_weights[531][6] = 4;
        layer_1_weights[532][6] = 0;
        layer_1_weights[533][6] = -1;
        layer_1_weights[534][6] = 1;
        layer_1_weights[535][6] = -2;
        layer_1_weights[536][6] = 0;
        layer_1_weights[537][6] = 2;
        layer_1_weights[538][6] = 2;
        layer_1_weights[539][6] = 2;
        layer_1_weights[540][6] = 1;
        layer_1_weights[541][6] = 0;
        layer_1_weights[542][6] = 1;
        layer_1_weights[543][6] = 2;
        layer_1_weights[544][6] = 1;
        layer_1_weights[545][6] = 3;
        layer_1_weights[546][6] = 2;
        layer_1_weights[547][6] = 1;
        layer_1_weights[548][6] = 0;
        layer_1_weights[549][6] = 0;
        layer_1_weights[550][6] = 1;
        layer_1_weights[551][6] = 0;
        layer_1_weights[552][6] = -2;
        layer_1_weights[553][6] = 0;
        layer_1_weights[554][6] = 1;
        layer_1_weights[555][6] = 1;
        layer_1_weights[556][6] = 3;
        layer_1_weights[557][6] = 5;
        layer_1_weights[558][6] = 2;
        layer_1_weights[559][6] = 2;
        layer_1_weights[560][6] = 1;
        layer_1_weights[561][6] = -1;
        layer_1_weights[562][6] = 3;
        layer_1_weights[563][6] = 1;
        layer_1_weights[564][6] = 2;
        layer_1_weights[565][6] = 1;
        layer_1_weights[566][6] = 1;
        layer_1_weights[567][6] = 0;
        layer_1_weights[568][6] = 2;
        layer_1_weights[569][6] = 1;
        layer_1_weights[570][6] = -1;
        layer_1_weights[571][6] = 1;
        layer_1_weights[572][6] = -1;
        layer_1_weights[573][6] = 0;
        layer_1_weights[574][6] = -1;
        layer_1_weights[575][6] = 0;
        layer_1_weights[576][6] = 2;
        layer_1_weights[577][6] = 2;
        layer_1_weights[578][6] = 1;
        layer_1_weights[579][6] = 1;
        layer_1_weights[580][6] = 2;
        layer_1_weights[581][6] = 0;
        layer_1_weights[582][6] = 0;
        layer_1_weights[583][6] = 1;
        layer_1_weights[584][6] = 5;
        layer_1_weights[585][6] = 3;
        layer_1_weights[586][6] = 1;
        layer_1_weights[587][6] = 3;
        layer_1_weights[588][6] = 0;
        layer_1_weights[589][6] = -1;
        layer_1_weights[590][6] = 0;
        layer_1_weights[591][6] = 1;
        layer_1_weights[592][6] = 1;
        layer_1_weights[593][6] = 3;
        layer_1_weights[594][6] = 1;
        layer_1_weights[595][6] = 1;
        layer_1_weights[596][6] = -1;
        layer_1_weights[597][6] = 0;
        layer_1_weights[598][6] = 0;
        layer_1_weights[599][6] = 0;
        layer_1_weights[600][6] = -2;
        layer_1_weights[601][6] = -2;
        layer_1_weights[602][6] = -1;
        layer_1_weights[603][6] = -1;
        layer_1_weights[604][6] = -1;
        layer_1_weights[605][6] = 0;
        layer_1_weights[606][6] = -1;
        layer_1_weights[607][6] = 0;
        layer_1_weights[608][6] = 0;
        layer_1_weights[609][6] = 0;
        layer_1_weights[610][6] = 2;
        layer_1_weights[611][6] = 0;
        layer_1_weights[612][6] = 5;
        layer_1_weights[613][6] = 3;
        layer_1_weights[614][6] = -2;
        layer_1_weights[615][6] = -1;
        layer_1_weights[616][6] = 1;
        layer_1_weights[617][6] = -2;
        layer_1_weights[618][6] = 0;
        layer_1_weights[619][6] = 2;
        layer_1_weights[620][6] = 1;
        layer_1_weights[621][6] = 0;
        layer_1_weights[622][6] = 1;
        layer_1_weights[623][6] = 0;
        layer_1_weights[624][6] = 0;
        layer_1_weights[625][6] = 0;
        layer_1_weights[626][6] = -1;
        layer_1_weights[627][6] = -2;
        layer_1_weights[628][6] = -1;
        layer_1_weights[629][6] = -1;
        layer_1_weights[630][6] = -1;
        layer_1_weights[631][6] = -1;
        layer_1_weights[632][6] = -1;
        layer_1_weights[633][6] = -1;
        layer_1_weights[634][6] = 0;
        layer_1_weights[635][6] = 0;
        layer_1_weights[636][6] = 0;
        layer_1_weights[637][6] = 1;
        layer_1_weights[638][6] = 2;
        layer_1_weights[639][6] = 3;
        layer_1_weights[640][6] = 7;
        layer_1_weights[641][6] = 6;
        layer_1_weights[642][6] = -2;
        layer_1_weights[643][6] = 0;
        layer_1_weights[644][6] = 0;
        layer_1_weights[645][6] = 0;
        layer_1_weights[646][6] = 1;
        layer_1_weights[647][6] = -1;
        layer_1_weights[648][6] = 1;
        layer_1_weights[649][6] = 1;
        layer_1_weights[650][6] = -1;
        layer_1_weights[651][6] = -1;
        layer_1_weights[652][6] = 1;
        layer_1_weights[653][6] = 1;
        layer_1_weights[654][6] = 1;
        layer_1_weights[655][6] = 2;
        layer_1_weights[656][6] = 0;
        layer_1_weights[657][6] = -1;
        layer_1_weights[658][6] = 0;
        layer_1_weights[659][6] = -1;
        layer_1_weights[660][6] = 0;
        layer_1_weights[661][6] = -1;
        layer_1_weights[662][6] = -2;
        layer_1_weights[663][6] = -1;
        layer_1_weights[664][6] = 1;
        layer_1_weights[665][6] = 0;
        layer_1_weights[666][6] = 1;
        layer_1_weights[667][6] = 3;
        layer_1_weights[668][6] = 3;
        layer_1_weights[669][6] = 4;
        layer_1_weights[670][6] = 3;
        layer_1_weights[671][6] = -1;
        layer_1_weights[672][6] = 0;
        layer_1_weights[673][6] = 0;
        layer_1_weights[674][6] = -1;
        layer_1_weights[675][6] = -3;
        layer_1_weights[676][6] = -2;
        layer_1_weights[677][6] = -1;
        layer_1_weights[678][6] = -2;
        layer_1_weights[679][6] = -1;
        layer_1_weights[680][6] = 0;
        layer_1_weights[681][6] = -2;
        layer_1_weights[682][6] = 1;
        layer_1_weights[683][6] = -1;
        layer_1_weights[684][6] = 0;
        layer_1_weights[685][6] = 0;
        layer_1_weights[686][6] = 0;
        layer_1_weights[687][6] = 1;
        layer_1_weights[688][6] = -1;
        layer_1_weights[689][6] = 1;
        layer_1_weights[690][6] = 1;
        layer_1_weights[691][6] = 2;
        layer_1_weights[692][6] = 1;
        layer_1_weights[693][6] = 3;
        layer_1_weights[694][6] = 3;
        layer_1_weights[695][6] = 4;
        layer_1_weights[696][6] = 8;
        layer_1_weights[697][6] = 3;
        layer_1_weights[698][6] = 2;
        layer_1_weights[699][6] = 0;
        layer_1_weights[700][6] = 0;
        layer_1_weights[701][6] = 0;
        layer_1_weights[702][6] = 3;
        layer_1_weights[703][6] = -2;
        layer_1_weights[704][6] = -2;
        layer_1_weights[705][6] = 0;
        layer_1_weights[706][6] = -3;
        layer_1_weights[707][6] = -1;
        layer_1_weights[708][6] = -2;
        layer_1_weights[709][6] = -2;
        layer_1_weights[710][6] = -3;
        layer_1_weights[711][6] = -2;
        layer_1_weights[712][6] = 1;
        layer_1_weights[713][6] = 1;
        layer_1_weights[714][6] = 0;
        layer_1_weights[715][6] = 1;
        layer_1_weights[716][6] = 2;
        layer_1_weights[717][6] = 2;
        layer_1_weights[718][6] = 3;
        layer_1_weights[719][6] = 1;
        layer_1_weights[720][6] = 4;
        layer_1_weights[721][6] = 4;
        layer_1_weights[722][6] = 4;
        layer_1_weights[723][6] = 1;
        layer_1_weights[724][6] = 4;
        layer_1_weights[725][6] = 2;
        layer_1_weights[726][6] = 1;
        layer_1_weights[727][6] = 0;
        layer_1_weights[728][6] = 1;
        layer_1_weights[729][6] = 0;
        layer_1_weights[730][6] = 0;
        layer_1_weights[731][6] = 2;
        layer_1_weights[732][6] = 0;
        layer_1_weights[733][6] = 2;
        layer_1_weights[734][6] = 3;
        layer_1_weights[735][6] = -3;
        layer_1_weights[736][6] = 0;
        layer_1_weights[737][6] = 1;
        layer_1_weights[738][6] = 2;
        layer_1_weights[739][6] = 3;
        layer_1_weights[740][6] = 1;
        layer_1_weights[741][6] = 1;
        layer_1_weights[742][6] = 2;
        layer_1_weights[743][6] = 3;
        layer_1_weights[744][6] = 0;
        layer_1_weights[745][6] = 1;
        layer_1_weights[746][6] = -1;
        layer_1_weights[747][6] = 1;
        layer_1_weights[748][6] = 3;
        layer_1_weights[749][6] = 3;
        layer_1_weights[750][6] = 2;
        layer_1_weights[751][6] = 1;
        layer_1_weights[752][6] = -1;
        layer_1_weights[753][6] = -2;
        layer_1_weights[754][6] = 0;
        layer_1_weights[755][6] = 1;
        layer_1_weights[756][6] = 0;
        layer_1_weights[757][6] = 1;
        layer_1_weights[758][6] = 1;
        layer_1_weights[759][6] = 0;
        layer_1_weights[760][6] = -2;
        layer_1_weights[761][6] = -4;
        layer_1_weights[762][6] = -3;
        layer_1_weights[763][6] = -6;
        layer_1_weights[764][6] = -5;
        layer_1_weights[765][6] = 1;
        layer_1_weights[766][6] = 1;
        layer_1_weights[767][6] = 2;
        layer_1_weights[768][6] = 1;
        layer_1_weights[769][6] = 0;
        layer_1_weights[770][6] = 2;
        layer_1_weights[771][6] = 1;
        layer_1_weights[772][6] = 0;
        layer_1_weights[773][6] = -2;
        layer_1_weights[774][6] = 1;
        layer_1_weights[775][6] = -1;
        layer_1_weights[776][6] = 0;
        layer_1_weights[777][6] = -2;
        layer_1_weights[778][6] = 0;
        layer_1_weights[779][6] = -3;
        layer_1_weights[780][6] = 0;
        layer_1_weights[781][6] = 0;
        layer_1_weights[782][6] = 0;
        layer_1_weights[783][6] = 0;
        layer_1_weights[0][7] = 1;
        layer_1_weights[1][7] = 0;
        layer_1_weights[2][7] = 0;
        layer_1_weights[3][7] = -1;
        layer_1_weights[4][7] = 0;
        layer_1_weights[5][7] = 0;
        layer_1_weights[6][7] = -1;
        layer_1_weights[7][7] = 0;
        layer_1_weights[8][7] = 0;
        layer_1_weights[9][7] = 0;
        layer_1_weights[10][7] = 0;
        layer_1_weights[11][7] = 0;
        layer_1_weights[12][7] = 0;
        layer_1_weights[13][7] = 2;
        layer_1_weights[14][7] = 3;
        layer_1_weights[15][7] = 0;
        layer_1_weights[16][7] = 0;
        layer_1_weights[17][7] = 0;
        layer_1_weights[18][7] = 1;
        layer_1_weights[19][7] = 0;
        layer_1_weights[20][7] = 0;
        layer_1_weights[21][7] = 0;
        layer_1_weights[22][7] = 0;
        layer_1_weights[23][7] = 0;
        layer_1_weights[24][7] = 0;
        layer_1_weights[25][7] = 0;
        layer_1_weights[26][7] = 0;
        layer_1_weights[27][7] = 0;
        layer_1_weights[28][7] = 0;
        layer_1_weights[29][7] = 0;
        layer_1_weights[30][7] = 0;
        layer_1_weights[31][7] = 1;
        layer_1_weights[32][7] = 0;
        layer_1_weights[33][7] = 0;
        layer_1_weights[34][7] = 0;
        layer_1_weights[35][7] = 0;
        layer_1_weights[36][7] = 3;
        layer_1_weights[37][7] = 2;
        layer_1_weights[38][7] = 2;
        layer_1_weights[39][7] = 3;
        layer_1_weights[40][7] = 0;
        layer_1_weights[41][7] = 3;
        layer_1_weights[42][7] = 4;
        layer_1_weights[43][7] = 3;
        layer_1_weights[44][7] = 4;
        layer_1_weights[45][7] = 2;
        layer_1_weights[46][7] = 3;
        layer_1_weights[47][7] = 2;
        layer_1_weights[48][7] = 2;
        layer_1_weights[49][7] = 0;
        layer_1_weights[50][7] = 1;
        layer_1_weights[51][7] = 0;
        layer_1_weights[52][7] = 0;
        layer_1_weights[53][7] = 0;
        layer_1_weights[54][7] = 0;
        layer_1_weights[55][7] = 0;
        layer_1_weights[56][7] = 0;
        layer_1_weights[57][7] = 0;
        layer_1_weights[58][7] = 2;
        layer_1_weights[59][7] = 0;
        layer_1_weights[60][7] = 2;
        layer_1_weights[61][7] = 0;
        layer_1_weights[62][7] = 1;
        layer_1_weights[63][7] = 0;
        layer_1_weights[64][7] = 1;
        layer_1_weights[65][7] = 3;
        layer_1_weights[66][7] = 1;
        layer_1_weights[67][7] = 1;
        layer_1_weights[68][7] = 2;
        layer_1_weights[69][7] = 2;
        layer_1_weights[70][7] = 3;
        layer_1_weights[71][7] = 1;
        layer_1_weights[72][7] = 2;
        layer_1_weights[73][7] = -4;
        layer_1_weights[74][7] = -1;
        layer_1_weights[75][7] = 0;
        layer_1_weights[76][7] = 1;
        layer_1_weights[77][7] = 2;
        layer_1_weights[78][7] = 0;
        layer_1_weights[79][7] = 1;
        layer_1_weights[80][7] = 3;
        layer_1_weights[81][7] = 3;
        layer_1_weights[82][7] = 0;
        layer_1_weights[83][7] = 0;
        layer_1_weights[84][7] = 0;
        layer_1_weights[85][7] = 1;
        layer_1_weights[86][7] = 2;
        layer_1_weights[87][7] = 2;
        layer_1_weights[88][7] = 0;
        layer_1_weights[89][7] = 2;
        layer_1_weights[90][7] = 1;
        layer_1_weights[91][7] = 0;
        layer_1_weights[92][7] = 3;
        layer_1_weights[93][7] = 4;
        layer_1_weights[94][7] = 2;
        layer_1_weights[95][7] = 3;
        layer_1_weights[96][7] = 4;
        layer_1_weights[97][7] = 1;
        layer_1_weights[98][7] = 2;
        layer_1_weights[99][7] = 3;
        layer_1_weights[100][7] = 2;
        layer_1_weights[101][7] = 2;
        layer_1_weights[102][7] = -1;
        layer_1_weights[103][7] = -2;
        layer_1_weights[104][7] = 3;
        layer_1_weights[105][7] = -1;
        layer_1_weights[106][7] = -3;
        layer_1_weights[107][7] = -7;
        layer_1_weights[108][7] = -2;
        layer_1_weights[109][7] = -1;
        layer_1_weights[110][7] = 0;
        layer_1_weights[111][7] = -1;
        layer_1_weights[112][7] = 0;
        layer_1_weights[113][7] = 2;
        layer_1_weights[114][7] = 4;
        layer_1_weights[115][7] = 2;
        layer_1_weights[116][7] = 5;
        layer_1_weights[117][7] = 1;
        layer_1_weights[118][7] = 0;
        layer_1_weights[119][7] = 2;
        layer_1_weights[120][7] = 2;
        layer_1_weights[121][7] = 0;
        layer_1_weights[122][7] = 1;
        layer_1_weights[123][7] = 3;
        layer_1_weights[124][7] = 3;
        layer_1_weights[125][7] = 2;
        layer_1_weights[126][7] = 3;
        layer_1_weights[127][7] = 3;
        layer_1_weights[128][7] = 4;
        layer_1_weights[129][7] = 1;
        layer_1_weights[130][7] = 2;
        layer_1_weights[131][7] = 0;
        layer_1_weights[132][7] = -2;
        layer_1_weights[133][7] = -1;
        layer_1_weights[134][7] = -1;
        layer_1_weights[135][7] = -5;
        layer_1_weights[136][7] = -5;
        layer_1_weights[137][7] = -4;
        layer_1_weights[138][7] = 3;
        layer_1_weights[139][7] = -1;
        layer_1_weights[140][7] = -1;
        layer_1_weights[141][7] = 1;
        layer_1_weights[142][7] = 1;
        layer_1_weights[143][7] = 2;
        layer_1_weights[144][7] = 3;
        layer_1_weights[145][7] = 1;
        layer_1_weights[146][7] = 0;
        layer_1_weights[147][7] = 0;
        layer_1_weights[148][7] = 1;
        layer_1_weights[149][7] = 2;
        layer_1_weights[150][7] = 1;
        layer_1_weights[151][7] = 0;
        layer_1_weights[152][7] = 1;
        layer_1_weights[153][7] = 2;
        layer_1_weights[154][7] = 2;
        layer_1_weights[155][7] = 2;
        layer_1_weights[156][7] = 0;
        layer_1_weights[157][7] = 0;
        layer_1_weights[158][7] = -1;
        layer_1_weights[159][7] = 0;
        layer_1_weights[160][7] = -2;
        layer_1_weights[161][7] = -1;
        layer_1_weights[162][7] = -1;
        layer_1_weights[163][7] = -1;
        layer_1_weights[164][7] = -2;
        layer_1_weights[165][7] = -3;
        layer_1_weights[166][7] = -2;
        layer_1_weights[167][7] = -2;
        layer_1_weights[168][7] = 0;
        layer_1_weights[169][7] = 0;
        layer_1_weights[170][7] = 1;
        layer_1_weights[171][7] = 4;
        layer_1_weights[172][7] = 2;
        layer_1_weights[173][7] = 1;
        layer_1_weights[174][7] = 0;
        layer_1_weights[175][7] = 1;
        layer_1_weights[176][7] = 0;
        layer_1_weights[177][7] = 0;
        layer_1_weights[178][7] = 1;
        layer_1_weights[179][7] = 1;
        layer_1_weights[180][7] = 0;
        layer_1_weights[181][7] = 0;
        layer_1_weights[182][7] = 0;
        layer_1_weights[183][7] = -1;
        layer_1_weights[184][7] = 0;
        layer_1_weights[185][7] = 0;
        layer_1_weights[186][7] = 1;
        layer_1_weights[187][7] = 1;
        layer_1_weights[188][7] = -1;
        layer_1_weights[189][7] = 1;
        layer_1_weights[190][7] = 1;
        layer_1_weights[191][7] = 0;
        layer_1_weights[192][7] = -3;
        layer_1_weights[193][7] = -3;
        layer_1_weights[194][7] = 1;
        layer_1_weights[195][7] = -2;
        layer_1_weights[196][7] = 0;
        layer_1_weights[197][7] = 6;
        layer_1_weights[198][7] = 2;
        layer_1_weights[199][7] = 2;
        layer_1_weights[200][7] = 2;
        layer_1_weights[201][7] = 0;
        layer_1_weights[202][7] = 0;
        layer_1_weights[203][7] = 0;
        layer_1_weights[204][7] = 0;
        layer_1_weights[205][7] = 2;
        layer_1_weights[206][7] = -1;
        layer_1_weights[207][7] = -1;
        layer_1_weights[208][7] = 0;
        layer_1_weights[209][7] = -1;
        layer_1_weights[210][7] = 1;
        layer_1_weights[211][7] = 1;
        layer_1_weights[212][7] = 2;
        layer_1_weights[213][7] = 2;
        layer_1_weights[214][7] = 2;
        layer_1_weights[215][7] = 1;
        layer_1_weights[216][7] = 1;
        layer_1_weights[217][7] = -1;
        layer_1_weights[218][7] = 0;
        layer_1_weights[219][7] = -1;
        layer_1_weights[220][7] = -3;
        layer_1_weights[221][7] = 0;
        layer_1_weights[222][7] = 1;
        layer_1_weights[223][7] = -2;
        layer_1_weights[224][7] = 3;
        layer_1_weights[225][7] = 5;
        layer_1_weights[226][7] = -2;
        layer_1_weights[227][7] = 2;
        layer_1_weights[228][7] = -1;
        layer_1_weights[229][7] = 0;
        layer_1_weights[230][7] = 3;
        layer_1_weights[231][7] = -1;
        layer_1_weights[232][7] = -3;
        layer_1_weights[233][7] = -2;
        layer_1_weights[234][7] = -4;
        layer_1_weights[235][7] = -5;
        layer_1_weights[236][7] = -3;
        layer_1_weights[237][7] = -2;
        layer_1_weights[238][7] = 0;
        layer_1_weights[239][7] = 3;
        layer_1_weights[240][7] = 3;
        layer_1_weights[241][7] = 3;
        layer_1_weights[242][7] = 2;
        layer_1_weights[243][7] = 2;
        layer_1_weights[244][7] = 1;
        layer_1_weights[245][7] = 1;
        layer_1_weights[246][7] = 2;
        layer_1_weights[247][7] = 0;
        layer_1_weights[248][7] = -1;
        layer_1_weights[249][7] = 1;
        layer_1_weights[250][7] = 1;
        layer_1_weights[251][7] = 3;
        layer_1_weights[252][7] = 2;
        layer_1_weights[253][7] = 3;
        layer_1_weights[254][7] = 0;
        layer_1_weights[255][7] = 2;
        layer_1_weights[256][7] = -4;
        layer_1_weights[257][7] = -4;
        layer_1_weights[258][7] = -3;
        layer_1_weights[259][7] = -7;
        layer_1_weights[260][7] = -4;
        layer_1_weights[261][7] = -5;
        layer_1_weights[262][7] = -3;
        layer_1_weights[263][7] = -4;
        layer_1_weights[264][7] = -5;
        layer_1_weights[265][7] = -2;
        layer_1_weights[266][7] = -1;
        layer_1_weights[267][7] = 1;
        layer_1_weights[268][7] = 3;
        layer_1_weights[269][7] = 2;
        layer_1_weights[270][7] = 2;
        layer_1_weights[271][7] = 1;
        layer_1_weights[272][7] = 2;
        layer_1_weights[273][7] = 0;
        layer_1_weights[274][7] = 0;
        layer_1_weights[275][7] = 1;
        layer_1_weights[276][7] = -2;
        layer_1_weights[277][7] = 0;
        layer_1_weights[278][7] = -4;
        layer_1_weights[279][7] = 1;
        layer_1_weights[280][7] = 1;
        layer_1_weights[281][7] = 3;
        layer_1_weights[282][7] = 3;
        layer_1_weights[283][7] = 0;
        layer_1_weights[284][7] = -4;
        layer_1_weights[285][7] = -7;
        layer_1_weights[286][7] = -6;
        layer_1_weights[287][7] = -6;
        layer_1_weights[288][7] = -4;
        layer_1_weights[289][7] = -4;
        layer_1_weights[290][7] = -3;
        layer_1_weights[291][7] = -2;
        layer_1_weights[292][7] = -4;
        layer_1_weights[293][7] = -3;
        layer_1_weights[294][7] = 0;
        layer_1_weights[295][7] = 1;
        layer_1_weights[296][7] = 1;
        layer_1_weights[297][7] = 1;
        layer_1_weights[298][7] = 0;
        layer_1_weights[299][7] = 1;
        layer_1_weights[300][7] = 0;
        layer_1_weights[301][7] = 0;
        layer_1_weights[302][7] = 3;
        layer_1_weights[303][7] = 0;
        layer_1_weights[304][7] = -4;
        layer_1_weights[305][7] = -2;
        layer_1_weights[306][7] = -1;
        layer_1_weights[307][7] = 2;
        layer_1_weights[308][7] = -1;
        layer_1_weights[309][7] = 3;
        layer_1_weights[310][7] = 1;
        layer_1_weights[311][7] = -4;
        layer_1_weights[312][7] = -5;
        layer_1_weights[313][7] = -5;
        layer_1_weights[314][7] = -4;
        layer_1_weights[315][7] = -2;
        layer_1_weights[316][7] = -2;
        layer_1_weights[317][7] = -1;
        layer_1_weights[318][7] = -1;
        layer_1_weights[319][7] = 1;
        layer_1_weights[320][7] = 0;
        layer_1_weights[321][7] = 1;
        layer_1_weights[322][7] = 1;
        layer_1_weights[323][7] = -1;
        layer_1_weights[324][7] = -2;
        layer_1_weights[325][7] = -1;
        layer_1_weights[326][7] = 0;
        layer_1_weights[327][7] = 1;
        layer_1_weights[328][7] = 1;
        layer_1_weights[329][7] = 1;
        layer_1_weights[330][7] = 1;
        layer_1_weights[331][7] = 1;
        layer_1_weights[332][7] = -2;
        layer_1_weights[333][7] = -3;
        layer_1_weights[334][7] = -3;
        layer_1_weights[335][7] = 3;
        layer_1_weights[336][7] = 0;
        layer_1_weights[337][7] = 1;
        layer_1_weights[338][7] = -1;
        layer_1_weights[339][7] = -1;
        layer_1_weights[340][7] = -3;
        layer_1_weights[341][7] = 0;
        layer_1_weights[342][7] = 0;
        layer_1_weights[343][7] = 2;
        layer_1_weights[344][7] = 0;
        layer_1_weights[345][7] = 2;
        layer_1_weights[346][7] = 2;
        layer_1_weights[347][7] = 2;
        layer_1_weights[348][7] = 1;
        layer_1_weights[349][7] = 0;
        layer_1_weights[350][7] = -1;
        layer_1_weights[351][7] = 1;
        layer_1_weights[352][7] = -1;
        layer_1_weights[353][7] = -1;
        layer_1_weights[354][7] = 1;
        layer_1_weights[355][7] = 0;
        layer_1_weights[356][7] = -1;
        layer_1_weights[357][7] = 0;
        layer_1_weights[358][7] = 0;
        layer_1_weights[359][7] = 1;
        layer_1_weights[360][7] = -2;
        layer_1_weights[361][7] = 0;
        layer_1_weights[362][7] = -3;
        layer_1_weights[363][7] = 2;
        layer_1_weights[364][7] = 0;
        layer_1_weights[365][7] = 1;
        layer_1_weights[366][7] = -1;
        layer_1_weights[367][7] = 0;
        layer_1_weights[368][7] = 1;
        layer_1_weights[369][7] = 1;
        layer_1_weights[370][7] = 0;
        layer_1_weights[371][7] = 3;
        layer_1_weights[372][7] = 2;
        layer_1_weights[373][7] = 3;
        layer_1_weights[374][7] = 2;
        layer_1_weights[375][7] = 1;
        layer_1_weights[376][7] = 1;
        layer_1_weights[377][7] = -1;
        layer_1_weights[378][7] = 0;
        layer_1_weights[379][7] = 0;
        layer_1_weights[380][7] = 0;
        layer_1_weights[381][7] = 0;
        layer_1_weights[382][7] = -1;
        layer_1_weights[383][7] = 0;
        layer_1_weights[384][7] = -2;
        layer_1_weights[385][7] = 1;
        layer_1_weights[386][7] = 0;
        layer_1_weights[387][7] = -1;
        layer_1_weights[388][7] = -1;
        layer_1_weights[389][7] = -1;
        layer_1_weights[390][7] = -2;
        layer_1_weights[391][7] = -1;
        layer_1_weights[392][7] = -2;
        layer_1_weights[393][7] = 1;
        layer_1_weights[394][7] = 3;
        layer_1_weights[395][7] = 2;
        layer_1_weights[396][7] = 1;
        layer_1_weights[397][7] = 4;
        layer_1_weights[398][7] = 3;
        layer_1_weights[399][7] = 0;
        layer_1_weights[400][7] = 4;
        layer_1_weights[401][7] = 2;
        layer_1_weights[402][7] = 1;
        layer_1_weights[403][7] = 1;
        layer_1_weights[404][7] = 0;
        layer_1_weights[405][7] = 1;
        layer_1_weights[406][7] = -1;
        layer_1_weights[407][7] = -1;
        layer_1_weights[408][7] = -1;
        layer_1_weights[409][7] = 0;
        layer_1_weights[410][7] = 0;
        layer_1_weights[411][7] = 0;
        layer_1_weights[412][7] = 0;
        layer_1_weights[413][7] = 0;
        layer_1_weights[414][7] = 0;
        layer_1_weights[415][7] = 0;
        layer_1_weights[416][7] = 1;
        layer_1_weights[417][7] = -3;
        layer_1_weights[418][7] = 2;
        layer_1_weights[419][7] = -1;
        layer_1_weights[420][7] = -2;
        layer_1_weights[421][7] = 1;
        layer_1_weights[422][7] = -1;
        layer_1_weights[423][7] = 1;
        layer_1_weights[424][7] = 2;
        layer_1_weights[425][7] = 4;
        layer_1_weights[426][7] = 1;
        layer_1_weights[427][7] = 1;
        layer_1_weights[428][7] = 0;
        layer_1_weights[429][7] = 0;
        layer_1_weights[430][7] = -2;
        layer_1_weights[431][7] = 0;
        layer_1_weights[432][7] = -2;
        layer_1_weights[433][7] = -1;
        layer_1_weights[434][7] = -1;
        layer_1_weights[435][7] = -1;
        layer_1_weights[436][7] = -1;
        layer_1_weights[437][7] = -1;
        layer_1_weights[438][7] = 0;
        layer_1_weights[439][7] = 0;
        layer_1_weights[440][7] = -2;
        layer_1_weights[441][7] = 1;
        layer_1_weights[442][7] = -1;
        layer_1_weights[443][7] = 1;
        layer_1_weights[444][7] = 3;
        layer_1_weights[445][7] = -4;
        layer_1_weights[446][7] = 3;
        layer_1_weights[447][7] = 1;
        layer_1_weights[448][7] = 0;
        layer_1_weights[449][7] = 3;
        layer_1_weights[450][7] = -1;
        layer_1_weights[451][7] = 2;
        layer_1_weights[452][7] = 2;
        layer_1_weights[453][7] = 2;
        layer_1_weights[454][7] = -1;
        layer_1_weights[455][7] = 0;
        layer_1_weights[456][7] = 1;
        layer_1_weights[457][7] = 1;
        layer_1_weights[458][7] = -1;
        layer_1_weights[459][7] = -1;
        layer_1_weights[460][7] = 0;
        layer_1_weights[461][7] = -2;
        layer_1_weights[462][7] = -1;
        layer_1_weights[463][7] = -1;
        layer_1_weights[464][7] = 0;
        layer_1_weights[465][7] = 1;
        layer_1_weights[466][7] = -1;
        layer_1_weights[467][7] = 0;
        layer_1_weights[468][7] = 0;
        layer_1_weights[469][7] = -2;
        layer_1_weights[470][7] = -2;
        layer_1_weights[471][7] = 0;
        layer_1_weights[472][7] = 1;
        layer_1_weights[473][7] = -4;
        layer_1_weights[474][7] = 1;
        layer_1_weights[475][7] = 1;
        layer_1_weights[476][7] = 0;
        layer_1_weights[477][7] = 3;
        layer_1_weights[478][7] = -1;
        layer_1_weights[479][7] = 0;
        layer_1_weights[480][7] = 0;
        layer_1_weights[481][7] = 2;
        layer_1_weights[482][7] = 0;
        layer_1_weights[483][7] = 0;
        layer_1_weights[484][7] = -1;
        layer_1_weights[485][7] = -2;
        layer_1_weights[486][7] = -1;
        layer_1_weights[487][7] = -2;
        layer_1_weights[488][7] = -2;
        layer_1_weights[489][7] = -1;
        layer_1_weights[490][7] = -3;
        layer_1_weights[491][7] = 0;
        layer_1_weights[492][7] = 0;
        layer_1_weights[493][7] = 1;
        layer_1_weights[494][7] = 0;
        layer_1_weights[495][7] = 0;
        layer_1_weights[496][7] = 0;
        layer_1_weights[497][7] = 0;
        layer_1_weights[498][7] = -1;
        layer_1_weights[499][7] = -3;
        layer_1_weights[500][7] = -2;
        layer_1_weights[501][7] = -1;
        layer_1_weights[502][7] = 0;
        layer_1_weights[503][7] = 3;
        layer_1_weights[504][7] = 2;
        layer_1_weights[505][7] = 1;
        layer_1_weights[506][7] = -1;
        layer_1_weights[507][7] = -2;
        layer_1_weights[508][7] = -1;
        layer_1_weights[509][7] = 0;
        layer_1_weights[510][7] = -1;
        layer_1_weights[511][7] = -1;
        layer_1_weights[512][7] = 0;
        layer_1_weights[513][7] = -1;
        layer_1_weights[514][7] = -1;
        layer_1_weights[515][7] = -2;
        layer_1_weights[516][7] = -2;
        layer_1_weights[517][7] = 0;
        layer_1_weights[518][7] = 1;
        layer_1_weights[519][7] = 1;
        layer_1_weights[520][7] = 0;
        layer_1_weights[521][7] = 1;
        layer_1_weights[522][7] = 1;
        layer_1_weights[523][7] = 0;
        layer_1_weights[524][7] = 0;
        layer_1_weights[525][7] = 1;
        layer_1_weights[526][7] = 0;
        layer_1_weights[527][7] = -1;
        layer_1_weights[528][7] = 0;
        layer_1_weights[529][7] = 2;
        layer_1_weights[530][7] = -1;
        layer_1_weights[531][7] = 3;
        layer_1_weights[532][7] = 0;
        layer_1_weights[533][7] = 4;
        layer_1_weights[534][7] = 1;
        layer_1_weights[535][7] = 0;
        layer_1_weights[536][7] = 0;
        layer_1_weights[537][7] = -1;
        layer_1_weights[538][7] = -2;
        layer_1_weights[539][7] = -1;
        layer_1_weights[540][7] = 0;
        layer_1_weights[541][7] = -1;
        layer_1_weights[542][7] = 0;
        layer_1_weights[543][7] = -1;
        layer_1_weights[544][7] = 0;
        layer_1_weights[545][7] = 2;
        layer_1_weights[546][7] = 1;
        layer_1_weights[547][7] = 1;
        layer_1_weights[548][7] = 0;
        layer_1_weights[549][7] = 2;
        layer_1_weights[550][7] = -1;
        layer_1_weights[551][7] = 0;
        layer_1_weights[552][7] = 0;
        layer_1_weights[553][7] = 0;
        layer_1_weights[554][7] = -2;
        layer_1_weights[555][7] = -1;
        layer_1_weights[556][7] = -1;
        layer_1_weights[557][7] = 0;
        layer_1_weights[558][7] = 1;
        layer_1_weights[559][7] = 3;
        layer_1_weights[560][7] = 0;
        layer_1_weights[561][7] = 3;
        layer_1_weights[562][7] = -3;
        layer_1_weights[563][7] = 0;
        layer_1_weights[564][7] = -1;
        layer_1_weights[565][7] = -2;
        layer_1_weights[566][7] = 0;
        layer_1_weights[567][7] = 0;
        layer_1_weights[568][7] = -1;
        layer_1_weights[569][7] = 1;
        layer_1_weights[570][7] = 1;
        layer_1_weights[571][7] = 2;
        layer_1_weights[572][7] = 2;
        layer_1_weights[573][7] = 2;
        layer_1_weights[574][7] = 1;
        layer_1_weights[575][7] = 1;
        layer_1_weights[576][7] = 0;
        layer_1_weights[577][7] = 0;
        layer_1_weights[578][7] = 2;
        layer_1_weights[579][7] = 0;
        layer_1_weights[580][7] = 1;
        layer_1_weights[581][7] = 1;
        layer_1_weights[582][7] = 0;
        layer_1_weights[583][7] = -3;
        layer_1_weights[584][7] = -3;
        layer_1_weights[585][7] = -1;
        layer_1_weights[586][7] = 1;
        layer_1_weights[587][7] = 3;
        layer_1_weights[588][7] = 0;
        layer_1_weights[589][7] = 1;
        layer_1_weights[590][7] = 4;
        layer_1_weights[591][7] = -1;
        layer_1_weights[592][7] = 0;
        layer_1_weights[593][7] = 0;
        layer_1_weights[594][7] = 0;
        layer_1_weights[595][7] = -1;
        layer_1_weights[596][7] = -1;
        layer_1_weights[597][7] = 1;
        layer_1_weights[598][7] = 0;
        layer_1_weights[599][7] = 0;
        layer_1_weights[600][7] = 1;
        layer_1_weights[601][7] = 1;
        layer_1_weights[602][7] = 1;
        layer_1_weights[603][7] = 0;
        layer_1_weights[604][7] = -1;
        layer_1_weights[605][7] = 0;
        layer_1_weights[606][7] = -1;
        layer_1_weights[607][7] = 0;
        layer_1_weights[608][7] = 0;
        layer_1_weights[609][7] = 1;
        layer_1_weights[610][7] = 0;
        layer_1_weights[611][7] = -2;
        layer_1_weights[612][7] = 0;
        layer_1_weights[613][7] = 2;
        layer_1_weights[614][7] = 3;
        layer_1_weights[615][7] = 1;
        layer_1_weights[616][7] = 0;
        layer_1_weights[617][7] = 1;
        layer_1_weights[618][7] = 2;
        layer_1_weights[619][7] = 2;
        layer_1_weights[620][7] = 0;
        layer_1_weights[621][7] = 1;
        layer_1_weights[622][7] = -1;
        layer_1_weights[623][7] = -1;
        layer_1_weights[624][7] = 2;
        layer_1_weights[625][7] = 0;
        layer_1_weights[626][7] = 0;
        layer_1_weights[627][7] = 0;
        layer_1_weights[628][7] = 0;
        layer_1_weights[629][7] = 1;
        layer_1_weights[630][7] = 0;
        layer_1_weights[631][7] = 1;
        layer_1_weights[632][7] = 0;
        layer_1_weights[633][7] = 2;
        layer_1_weights[634][7] = 1;
        layer_1_weights[635][7] = -2;
        layer_1_weights[636][7] = 1;
        layer_1_weights[637][7] = -2;
        layer_1_weights[638][7] = 0;
        layer_1_weights[639][7] = 2;
        layer_1_weights[640][7] = 0;
        layer_1_weights[641][7] = -2;
        layer_1_weights[642][7] = 2;
        layer_1_weights[643][7] = 2;
        layer_1_weights[644][7] = 0;
        layer_1_weights[645][7] = 1;
        layer_1_weights[646][7] = 3;
        layer_1_weights[647][7] = 1;
        layer_1_weights[648][7] = 1;
        layer_1_weights[649][7] = -1;
        layer_1_weights[650][7] = -1;
        layer_1_weights[651][7] = 0;
        layer_1_weights[652][7] = 0;
        layer_1_weights[653][7] = 1;
        layer_1_weights[654][7] = 2;
        layer_1_weights[655][7] = 1;
        layer_1_weights[656][7] = 2;
        layer_1_weights[657][7] = 1;
        layer_1_weights[658][7] = 2;
        layer_1_weights[659][7] = 0;
        layer_1_weights[660][7] = 1;
        layer_1_weights[661][7] = 0;
        layer_1_weights[662][7] = 0;
        layer_1_weights[663][7] = 1;
        layer_1_weights[664][7] = -2;
        layer_1_weights[665][7] = 2;
        layer_1_weights[666][7] = 0;
        layer_1_weights[667][7] = 2;
        layer_1_weights[668][7] = 3;
        layer_1_weights[669][7] = 3;
        layer_1_weights[670][7] = 3;
        layer_1_weights[671][7] = 0;
        layer_1_weights[672][7] = 0;
        layer_1_weights[673][7] = 0;
        layer_1_weights[674][7] = -2;
        layer_1_weights[675][7] = 3;
        layer_1_weights[676][7] = 1;
        layer_1_weights[677][7] = -2;
        layer_1_weights[678][7] = 0;
        layer_1_weights[679][7] = 0;
        layer_1_weights[680][7] = 1;
        layer_1_weights[681][7] = 0;
        layer_1_weights[682][7] = 2;
        layer_1_weights[683][7] = 0;
        layer_1_weights[684][7] = 1;
        layer_1_weights[685][7] = 1;
        layer_1_weights[686][7] = 0;
        layer_1_weights[687][7] = 2;
        layer_1_weights[688][7] = 1;
        layer_1_weights[689][7] = 1;
        layer_1_weights[690][7] = 0;
        layer_1_weights[691][7] = -2;
        layer_1_weights[692][7] = 0;
        layer_1_weights[693][7] = 2;
        layer_1_weights[694][7] = 2;
        layer_1_weights[695][7] = -2;
        layer_1_weights[696][7] = 0;
        layer_1_weights[697][7] = 1;
        layer_1_weights[698][7] = 1;
        layer_1_weights[699][7] = 1;
        layer_1_weights[700][7] = 0;
        layer_1_weights[701][7] = 0;
        layer_1_weights[702][7] = 0;
        layer_1_weights[703][7] = 1;
        layer_1_weights[704][7] = 2;
        layer_1_weights[705][7] = 1;
        layer_1_weights[706][7] = 1;
        layer_1_weights[707][7] = 3;
        layer_1_weights[708][7] = 3;
        layer_1_weights[709][7] = 1;
        layer_1_weights[710][7] = 2;
        layer_1_weights[711][7] = -1;
        layer_1_weights[712][7] = 0;
        layer_1_weights[713][7] = 1;
        layer_1_weights[714][7] = 0;
        layer_1_weights[715][7] = -1;
        layer_1_weights[716][7] = -1;
        layer_1_weights[717][7] = -4;
        layer_1_weights[718][7] = -3;
        layer_1_weights[719][7] = 0;
        layer_1_weights[720][7] = 2;
        layer_1_weights[721][7] = -2;
        layer_1_weights[722][7] = -3;
        layer_1_weights[723][7] = -2;
        layer_1_weights[724][7] = -1;
        layer_1_weights[725][7] = 0;
        layer_1_weights[726][7] = 0;
        layer_1_weights[727][7] = 0;
        layer_1_weights[728][7] = 0;
        layer_1_weights[729][7] = 0;
        layer_1_weights[730][7] = 0;
        layer_1_weights[731][7] = 1;
        layer_1_weights[732][7] = -1;
        layer_1_weights[733][7] = 1;
        layer_1_weights[734][7] = -2;
        layer_1_weights[735][7] = 0;
        layer_1_weights[736][7] = -2;
        layer_1_weights[737][7] = -1;
        layer_1_weights[738][7] = 0;
        layer_1_weights[739][7] = -2;
        layer_1_weights[740][7] = 1;
        layer_1_weights[741][7] = 2;
        layer_1_weights[742][7] = 1;
        layer_1_weights[743][7] = -1;
        layer_1_weights[744][7] = 0;
        layer_1_weights[745][7] = -3;
        layer_1_weights[746][7] = -2;
        layer_1_weights[747][7] = -1;
        layer_1_weights[748][7] = 0;
        layer_1_weights[749][7] = 2;
        layer_1_weights[750][7] = 1;
        layer_1_weights[751][7] = 1;
        layer_1_weights[752][7] = 1;
        layer_1_weights[753][7] = 2;
        layer_1_weights[754][7] = 0;
        layer_1_weights[755][7] = 0;
        layer_1_weights[756][7] = 0;
        layer_1_weights[757][7] = 1;
        layer_1_weights[758][7] = 0;
        layer_1_weights[759][7] = 0;
        layer_1_weights[760][7] = 0;
        layer_1_weights[761][7] = 1;
        layer_1_weights[762][7] = -1;
        layer_1_weights[763][7] = -1;
        layer_1_weights[764][7] = 0;
        layer_1_weights[765][7] = -2;
        layer_1_weights[766][7] = -1;
        layer_1_weights[767][7] = 0;
        layer_1_weights[768][7] = 0;
        layer_1_weights[769][7] = 2;
        layer_1_weights[770][7] = 3;
        layer_1_weights[771][7] = 3;
        layer_1_weights[772][7] = 3;
        layer_1_weights[773][7] = 1;
        layer_1_weights[774][7] = 0;
        layer_1_weights[775][7] = 3;
        layer_1_weights[776][7] = 0;
        layer_1_weights[777][7] = 0;
        layer_1_weights[778][7] = 0;
        layer_1_weights[779][7] = -1;
        layer_1_weights[780][7] = -1;
        layer_1_weights[781][7] = -1;
        layer_1_weights[782][7] = 0;
        layer_1_weights[783][7] = -1;
        layer_1_weights[0][8] = -1;
        layer_1_weights[1][8] = 0;
        layer_1_weights[2][8] = 0;
        layer_1_weights[3][8] = -1;
        layer_1_weights[4][8] = 0;
        layer_1_weights[5][8] = 0;
        layer_1_weights[6][8] = 0;
        layer_1_weights[7][8] = 0;
        layer_1_weights[8][8] = 1;
        layer_1_weights[9][8] = 0;
        layer_1_weights[10][8] = 0;
        layer_1_weights[11][8] = 0;
        layer_1_weights[12][8] = 2;
        layer_1_weights[13][8] = -2;
        layer_1_weights[14][8] = -2;
        layer_1_weights[15][8] = -1;
        layer_1_weights[16][8] = 0;
        layer_1_weights[17][8] = -1;
        layer_1_weights[18][8] = 1;
        layer_1_weights[19][8] = 0;
        layer_1_weights[20][8] = -1;
        layer_1_weights[21][8] = 0;
        layer_1_weights[22][8] = 0;
        layer_1_weights[23][8] = 0;
        layer_1_weights[24][8] = 0;
        layer_1_weights[25][8] = 0;
        layer_1_weights[26][8] = 1;
        layer_1_weights[27][8] = 0;
        layer_1_weights[28][8] = 0;
        layer_1_weights[29][8] = 0;
        layer_1_weights[30][8] = 0;
        layer_1_weights[31][8] = 0;
        layer_1_weights[32][8] = 0;
        layer_1_weights[33][8] = 2;
        layer_1_weights[34][8] = 4;
        layer_1_weights[35][8] = 5;
        layer_1_weights[36][8] = 3;
        layer_1_weights[37][8] = 2;
        layer_1_weights[38][8] = 3;
        layer_1_weights[39][8] = 2;
        layer_1_weights[40][8] = 3;
        layer_1_weights[41][8] = 3;
        layer_1_weights[42][8] = 2;
        layer_1_weights[43][8] = 1;
        layer_1_weights[44][8] = 1;
        layer_1_weights[45][8] = 3;
        layer_1_weights[46][8] = 1;
        layer_1_weights[47][8] = 4;
        layer_1_weights[48][8] = 5;
        layer_1_weights[49][8] = 3;
        layer_1_weights[50][8] = 2;
        layer_1_weights[51][8] = 1;
        layer_1_weights[52][8] = 0;
        layer_1_weights[53][8] = 0;
        layer_1_weights[54][8] = 0;
        layer_1_weights[55][8] = -1;
        layer_1_weights[56][8] = 1;
        layer_1_weights[57][8] = 0;
        layer_1_weights[58][8] = 1;
        layer_1_weights[59][8] = -1;
        layer_1_weights[60][8] = 2;
        layer_1_weights[61][8] = 0;
        layer_1_weights[62][8] = 5;
        layer_1_weights[63][8] = 4;
        layer_1_weights[64][8] = -1;
        layer_1_weights[65][8] = -1;
        layer_1_weights[66][8] = 0;
        layer_1_weights[67][8] = 4;
        layer_1_weights[68][8] = 0;
        layer_1_weights[69][8] = 0;
        layer_1_weights[70][8] = -3;
        layer_1_weights[71][8] = -1;
        layer_1_weights[72][8] = -3;
        layer_1_weights[73][8] = 1;
        layer_1_weights[74][8] = 0;
        layer_1_weights[75][8] = 1;
        layer_1_weights[76][8] = 0;
        layer_1_weights[77][8] = 2;
        layer_1_weights[78][8] = 6;
        layer_1_weights[79][8] = 2;
        layer_1_weights[80][8] = -1;
        layer_1_weights[81][8] = 0;
        layer_1_weights[82][8] = 0;
        layer_1_weights[83][8] = -1;
        layer_1_weights[84][8] = 0;
        layer_1_weights[85][8] = -1;
        layer_1_weights[86][8] = -2;
        layer_1_weights[87][8] = 3;
        layer_1_weights[88][8] = 4;
        layer_1_weights[89][8] = 2;
        layer_1_weights[90][8] = -1;
        layer_1_weights[91][8] = 2;
        layer_1_weights[92][8] = 1;
        layer_1_weights[93][8] = 1;
        layer_1_weights[94][8] = 2;
        layer_1_weights[95][8] = 5;
        layer_1_weights[96][8] = 2;
        layer_1_weights[97][8] = 2;
        layer_1_weights[98][8] = 2;
        layer_1_weights[99][8] = 2;
        layer_1_weights[100][8] = 1;
        layer_1_weights[101][8] = 0;
        layer_1_weights[102][8] = 1;
        layer_1_weights[103][8] = 1;
        layer_1_weights[104][8] = 2;
        layer_1_weights[105][8] = 2;
        layer_1_weights[106][8] = -2;
        layer_1_weights[107][8] = 0;
        layer_1_weights[108][8] = 3;
        layer_1_weights[109][8] = 2;
        layer_1_weights[110][8] = 3;
        layer_1_weights[111][8] = 0;
        layer_1_weights[112][8] = 0;
        layer_1_weights[113][8] = 2;
        layer_1_weights[114][8] = -1;
        layer_1_weights[115][8] = 1;
        layer_1_weights[116][8] = 0;
        layer_1_weights[117][8] = -1;
        layer_1_weights[118][8] = 1;
        layer_1_weights[119][8] = 2;
        layer_1_weights[120][8] = 2;
        layer_1_weights[121][8] = 2;
        layer_1_weights[122][8] = 3;
        layer_1_weights[123][8] = 1;
        layer_1_weights[124][8] = 0;
        layer_1_weights[125][8] = 1;
        layer_1_weights[126][8] = 1;
        layer_1_weights[127][8] = 1;
        layer_1_weights[128][8] = 2;
        layer_1_weights[129][8] = 2;
        layer_1_weights[130][8] = 1;
        layer_1_weights[131][8] = 3;
        layer_1_weights[132][8] = 1;
        layer_1_weights[133][8] = 1;
        layer_1_weights[134][8] = 2;
        layer_1_weights[135][8] = 1;
        layer_1_weights[136][8] = 2;
        layer_1_weights[137][8] = 4;
        layer_1_weights[138][8] = 0;
        layer_1_weights[139][8] = 2;
        layer_1_weights[140][8] = -1;
        layer_1_weights[141][8] = -1;
        layer_1_weights[142][8] = -1;
        layer_1_weights[143][8] = 3;
        layer_1_weights[144][8] = 1;
        layer_1_weights[145][8] = -1;
        layer_1_weights[146][8] = -1;
        layer_1_weights[147][8] = 1;
        layer_1_weights[148][8] = 1;
        layer_1_weights[149][8] = -1;
        layer_1_weights[150][8] = 2;
        layer_1_weights[151][8] = 0;
        layer_1_weights[152][8] = 0;
        layer_1_weights[153][8] = 0;
        layer_1_weights[154][8] = 0;
        layer_1_weights[155][8] = 0;
        layer_1_weights[156][8] = 0;
        layer_1_weights[157][8] = 1;
        layer_1_weights[158][8] = 1;
        layer_1_weights[159][8] = 2;
        layer_1_weights[160][8] = 2;
        layer_1_weights[161][8] = 2;
        layer_1_weights[162][8] = 1;
        layer_1_weights[163][8] = 3;
        layer_1_weights[164][8] = 3;
        layer_1_weights[165][8] = 0;
        layer_1_weights[166][8] = 3;
        layer_1_weights[167][8] = 3;
        layer_1_weights[168][8] = -1;
        layer_1_weights[169][8] = 0;
        layer_1_weights[170][8] = 0;
        layer_1_weights[171][8] = -2;
        layer_1_weights[172][8] = 1;
        layer_1_weights[173][8] = 0;
        layer_1_weights[174][8] = 1;
        layer_1_weights[175][8] = 1;
        layer_1_weights[176][8] = -1;
        layer_1_weights[177][8] = 0;
        layer_1_weights[178][8] = 0;
        layer_1_weights[179][8] = -1;
        layer_1_weights[180][8] = -1;
        layer_1_weights[181][8] = -1;
        layer_1_weights[182][8] = -1;
        layer_1_weights[183][8] = -1;
        layer_1_weights[184][8] = -1;
        layer_1_weights[185][8] = -2;
        layer_1_weights[186][8] = -2;
        layer_1_weights[187][8] = -2;
        layer_1_weights[188][8] = 0;
        layer_1_weights[189][8] = -1;
        layer_1_weights[190][8] = 2;
        layer_1_weights[191][8] = 3;
        layer_1_weights[192][8] = 5;
        layer_1_weights[193][8] = 3;
        layer_1_weights[194][8] = 4;
        layer_1_weights[195][8] = 1;
        layer_1_weights[196][8] = -1;
        layer_1_weights[197][8] = 2;
        layer_1_weights[198][8] = 0;
        layer_1_weights[199][8] = 1;
        layer_1_weights[200][8] = 3;
        layer_1_weights[201][8] = 5;
        layer_1_weights[202][8] = 1;
        layer_1_weights[203][8] = 1;
        layer_1_weights[204][8] = 1;
        layer_1_weights[205][8] = 1;
        layer_1_weights[206][8] = 0;
        layer_1_weights[207][8] = 0;
        layer_1_weights[208][8] = 0;
        layer_1_weights[209][8] = 0;
        layer_1_weights[210][8] = -1;
        layer_1_weights[211][8] = -1;
        layer_1_weights[212][8] = -1;
        layer_1_weights[213][8] = -1;
        layer_1_weights[214][8] = -2;
        layer_1_weights[215][8] = -2;
        layer_1_weights[216][8] = 0;
        layer_1_weights[217][8] = -1;
        layer_1_weights[218][8] = -1;
        layer_1_weights[219][8] = 2;
        layer_1_weights[220][8] = 3;
        layer_1_weights[221][8] = 2;
        layer_1_weights[222][8] = 7;
        layer_1_weights[223][8] = 1;
        layer_1_weights[224][8] = 3;
        layer_1_weights[225][8] = -2;
        layer_1_weights[226][8] = 0;
        layer_1_weights[227][8] = 0;
        layer_1_weights[228][8] = 0;
        layer_1_weights[229][8] = 1;
        layer_1_weights[230][8] = 0;
        layer_1_weights[231][8] = -1;
        layer_1_weights[232][8] = -1;
        layer_1_weights[233][8] = 1;
        layer_1_weights[234][8] = 0;
        layer_1_weights[235][8] = 0;
        layer_1_weights[236][8] = 0;
        layer_1_weights[237][8] = 0;
        layer_1_weights[238][8] = 0;
        layer_1_weights[239][8] = 0;
        layer_1_weights[240][8] = 1;
        layer_1_weights[241][8] = 0;
        layer_1_weights[242][8] = 1;
        layer_1_weights[243][8] = 1;
        layer_1_weights[244][8] = 1;
        layer_1_weights[245][8] = 1;
        layer_1_weights[246][8] = 1;
        layer_1_weights[247][8] = 3;
        layer_1_weights[248][8] = 2;
        layer_1_weights[249][8] = 3;
        layer_1_weights[250][8] = 3;
        layer_1_weights[251][8] = 1;
        layer_1_weights[252][8] = -2;
        layer_1_weights[253][8] = -5;
        layer_1_weights[254][8] = 3;
        layer_1_weights[255][8] = 0;
        layer_1_weights[256][8] = 3;
        layer_1_weights[257][8] = -1;
        layer_1_weights[258][8] = -1;
        layer_1_weights[259][8] = 1;
        layer_1_weights[260][8] = 1;
        layer_1_weights[261][8] = -2;
        layer_1_weights[262][8] = -1;
        layer_1_weights[263][8] = 0;
        layer_1_weights[264][8] = -1;
        layer_1_weights[265][8] = 0;
        layer_1_weights[266][8] = 0;
        layer_1_weights[267][8] = 0;
        layer_1_weights[268][8] = 1;
        layer_1_weights[269][8] = 1;
        layer_1_weights[270][8] = 0;
        layer_1_weights[271][8] = 0;
        layer_1_weights[272][8] = 1;
        layer_1_weights[273][8] = 0;
        layer_1_weights[274][8] = -1;
        layer_1_weights[275][8] = 2;
        layer_1_weights[276][8] = 1;
        layer_1_weights[277][8] = 2;
        layer_1_weights[278][8] = 0;
        layer_1_weights[279][8] = -2;
        layer_1_weights[280][8] = -1;
        layer_1_weights[281][8] = -5;
        layer_1_weights[282][8] = 1;
        layer_1_weights[283][8] = 0;
        layer_1_weights[284][8] = 2;
        layer_1_weights[285][8] = -2;
        layer_1_weights[286][8] = 0;
        layer_1_weights[287][8] = 1;
        layer_1_weights[288][8] = 1;
        layer_1_weights[289][8] = 0;
        layer_1_weights[290][8] = -2;
        layer_1_weights[291][8] = -1;
        layer_1_weights[292][8] = 0;
        layer_1_weights[293][8] = 0;
        layer_1_weights[294][8] = -1;
        layer_1_weights[295][8] = -1;
        layer_1_weights[296][8] = 0;
        layer_1_weights[297][8] = 0;
        layer_1_weights[298][8] = 1;
        layer_1_weights[299][8] = 1;
        layer_1_weights[300][8] = 1;
        layer_1_weights[301][8] = 0;
        layer_1_weights[302][8] = -1;
        layer_1_weights[303][8] = 0;
        layer_1_weights[304][8] = 4;
        layer_1_weights[305][8] = 1;
        layer_1_weights[306][8] = 0;
        layer_1_weights[307][8] = -5;
        layer_1_weights[308][8] = -2;
        layer_1_weights[309][8] = 1;
        layer_1_weights[310][8] = -2;
        layer_1_weights[311][8] = 3;
        layer_1_weights[312][8] = -2;
        layer_1_weights[313][8] = -1;
        layer_1_weights[314][8] = 1;
        layer_1_weights[315][8] = 0;
        layer_1_weights[316][8] = 0;
        layer_1_weights[317][8] = 0;
        layer_1_weights[318][8] = 0;
        layer_1_weights[319][8] = 0;
        layer_1_weights[320][8] = 1;
        layer_1_weights[321][8] = 2;
        layer_1_weights[322][8] = 0;
        layer_1_weights[323][8] = -1;
        layer_1_weights[324][8] = 0;
        layer_1_weights[325][8] = -1;
        layer_1_weights[326][8] = 0;
        layer_1_weights[327][8] = 0;
        layer_1_weights[328][8] = -1;
        layer_1_weights[329][8] = 0;
        layer_1_weights[330][8] = -3;
        layer_1_weights[331][8] = -1;
        layer_1_weights[332][8] = 2;
        layer_1_weights[333][8] = 0;
        layer_1_weights[334][8] = 1;
        layer_1_weights[335][8] = -1;
        layer_1_weights[336][8] = -1;
        layer_1_weights[337][8] = -5;
        layer_1_weights[338][8] = -4;
        layer_1_weights[339][8] = -1;
        layer_1_weights[340][8] = -2;
        layer_1_weights[341][8] = -1;
        layer_1_weights[342][8] = 1;
        layer_1_weights[343][8] = -1;
        layer_1_weights[344][8] = -1;
        layer_1_weights[345][8] = -2;
        layer_1_weights[346][8] = 1;
        layer_1_weights[347][8] = 1;
        layer_1_weights[348][8] = 2;
        layer_1_weights[349][8] = 2;
        layer_1_weights[350][8] = 0;
        layer_1_weights[351][8] = 1;
        layer_1_weights[352][8] = -1;
        layer_1_weights[353][8] = -1;
        layer_1_weights[354][8] = -1;
        layer_1_weights[355][8] = 0;
        layer_1_weights[356][8] = 0;
        layer_1_weights[357][8] = -2;
        layer_1_weights[358][8] = -2;
        layer_1_weights[359][8] = 0;
        layer_1_weights[360][8] = 2;
        layer_1_weights[361][8] = 1;
        layer_1_weights[362][8] = 2;
        layer_1_weights[363][8] = -2;
        layer_1_weights[364][8] = 0;
        layer_1_weights[365][8] = -1;
        layer_1_weights[366][8] = 0;
        layer_1_weights[367][8] = 1;
        layer_1_weights[368][8] = -2;
        layer_1_weights[369][8] = 0;
        layer_1_weights[370][8] = 0;
        layer_1_weights[371][8] = 0;
        layer_1_weights[372][8] = -1;
        layer_1_weights[373][8] = 1;
        layer_1_weights[374][8] = 1;
        layer_1_weights[375][8] = 1;
        layer_1_weights[376][8] = 2;
        layer_1_weights[377][8] = 3;
        layer_1_weights[378][8] = 0;
        layer_1_weights[379][8] = -1;
        layer_1_weights[380][8] = -1;
        layer_1_weights[381][8] = 0;
        layer_1_weights[382][8] = 1;
        layer_1_weights[383][8] = 2;
        layer_1_weights[384][8] = -1;
        layer_1_weights[385][8] = -1;
        layer_1_weights[386][8] = -1;
        layer_1_weights[387][8] = 1;
        layer_1_weights[388][8] = 0;
        layer_1_weights[389][8] = -1;
        layer_1_weights[390][8] = -2;
        layer_1_weights[391][8] = 1;
        layer_1_weights[392][8] = 3;
        layer_1_weights[393][8] = 1;
        layer_1_weights[394][8] = -4;
        layer_1_weights[395][8] = -2;
        layer_1_weights[396][8] = 1;
        layer_1_weights[397][8] = 0;
        layer_1_weights[398][8] = 0;
        layer_1_weights[399][8] = 1;
        layer_1_weights[400][8] = 1;
        layer_1_weights[401][8] = 0;
        layer_1_weights[402][8] = 2;
        layer_1_weights[403][8] = 2;
        layer_1_weights[404][8] = 3;
        layer_1_weights[405][8] = 2;
        layer_1_weights[406][8] = 0;
        layer_1_weights[407][8] = -1;
        layer_1_weights[408][8] = -1;
        layer_1_weights[409][8] = 0;
        layer_1_weights[410][8] = 0;
        layer_1_weights[411][8] = 0;
        layer_1_weights[412][8] = -1;
        layer_1_weights[413][8] = -1;
        layer_1_weights[414][8] = 0;
        layer_1_weights[415][8] = 3;
        layer_1_weights[416][8] = -1;
        layer_1_weights[417][8] = -1;
        layer_1_weights[418][8] = -3;
        layer_1_weights[419][8] = -3;
        layer_1_weights[420][8] = 2;
        layer_1_weights[421][8] = 1;
        layer_1_weights[422][8] = 3;
        layer_1_weights[423][8] = 2;
        layer_1_weights[424][8] = 1;
        layer_1_weights[425][8] = 0;
        layer_1_weights[426][8] = 0;
        layer_1_weights[427][8] = 1;
        layer_1_weights[428][8] = -1;
        layer_1_weights[429][8] = 0;
        layer_1_weights[430][8] = 0;
        layer_1_weights[431][8] = 2;
        layer_1_weights[432][8] = 2;
        layer_1_weights[433][8] = 2;
        layer_1_weights[434][8] = 1;
        layer_1_weights[435][8] = 1;
        layer_1_weights[436][8] = -1;
        layer_1_weights[437][8] = 1;
        layer_1_weights[438][8] = 0;
        layer_1_weights[439][8] = 1;
        layer_1_weights[440][8] = 1;
        layer_1_weights[441][8] = 0;
        layer_1_weights[442][8] = 2;
        layer_1_weights[443][8] = 1;
        layer_1_weights[444][8] = 2;
        layer_1_weights[445][8] = 3;
        layer_1_weights[446][8] = -3;
        layer_1_weights[447][8] = -3;
        layer_1_weights[448][8] = -2;
        layer_1_weights[449][8] = 3;
        layer_1_weights[450][8] = 0;
        layer_1_weights[451][8] = 1;
        layer_1_weights[452][8] = 0;
        layer_1_weights[453][8] = 1;
        layer_1_weights[454][8] = 0;
        layer_1_weights[455][8] = 2;
        layer_1_weights[456][8] = 0;
        layer_1_weights[457][8] = -1;
        layer_1_weights[458][8] = -1;
        layer_1_weights[459][8] = 1;
        layer_1_weights[460][8] = 2;
        layer_1_weights[461][8] = 1;
        layer_1_weights[462][8] = 0;
        layer_1_weights[463][8] = 0;
        layer_1_weights[464][8] = -1;
        layer_1_weights[465][8] = 1;
        layer_1_weights[466][8] = 1;
        layer_1_weights[467][8] = 2;
        layer_1_weights[468][8] = 2;
        layer_1_weights[469][8] = 0;
        layer_1_weights[470][8] = 0;
        layer_1_weights[471][8] = 0;
        layer_1_weights[472][8] = 2;
        layer_1_weights[473][8] = 2;
        layer_1_weights[474][8] = -4;
        layer_1_weights[475][8] = -2;
        layer_1_weights[476][8] = 0;
        layer_1_weights[477][8] = 2;
        layer_1_weights[478][8] = 1;
        layer_1_weights[479][8] = 3;
        layer_1_weights[480][8] = 2;
        layer_1_weights[481][8] = 1;
        layer_1_weights[482][8] = 1;
        layer_1_weights[483][8] = 0;
        layer_1_weights[484][8] = -2;
        layer_1_weights[485][8] = -1;
        layer_1_weights[486][8] = -1;
        layer_1_weights[487][8] = 0;
        layer_1_weights[488][8] = 1;
        layer_1_weights[489][8] = 0;
        layer_1_weights[490][8] = -3;
        layer_1_weights[491][8] = 0;
        layer_1_weights[492][8] = 0;
        layer_1_weights[493][8] = 2;
        layer_1_weights[494][8] = 1;
        layer_1_weights[495][8] = 1;
        layer_1_weights[496][8] = 1;
        layer_1_weights[497][8] = 2;
        layer_1_weights[498][8] = 0;
        layer_1_weights[499][8] = 4;
        layer_1_weights[500][8] = 2;
        layer_1_weights[501][8] = -1;
        layer_1_weights[502][8] = -4;
        layer_1_weights[503][8] = 0;
        layer_1_weights[504][8] = -3;
        layer_1_weights[505][8] = -1;
        layer_1_weights[506][8] = 0;
        layer_1_weights[507][8] = 3;
        layer_1_weights[508][8] = 2;
        layer_1_weights[509][8] = 4;
        layer_1_weights[510][8] = 1;
        layer_1_weights[511][8] = 0;
        layer_1_weights[512][8] = 0;
        layer_1_weights[513][8] = 0;
        layer_1_weights[514][8] = 0;
        layer_1_weights[515][8] = 1;
        layer_1_weights[516][8] = 1;
        layer_1_weights[517][8] = 1;
        layer_1_weights[518][8] = -1;
        layer_1_weights[519][8] = 1;
        layer_1_weights[520][8] = 2;
        layer_1_weights[521][8] = 2;
        layer_1_weights[522][8] = 1;
        layer_1_weights[523][8] = 0;
        layer_1_weights[524][8] = -1;
        layer_1_weights[525][8] = 1;
        layer_1_weights[526][8] = -2;
        layer_1_weights[527][8] = 2;
        layer_1_weights[528][8] = 1;
        layer_1_weights[529][8] = -1;
        layer_1_weights[530][8] = -5;
        layer_1_weights[531][8] = -4;
        layer_1_weights[532][8] = 0;
        layer_1_weights[533][8] = -2;
        layer_1_weights[534][8] = 0;
        layer_1_weights[535][8] = 2;
        layer_1_weights[536][8] = 2;
        layer_1_weights[537][8] = 3;
        layer_1_weights[538][8] = 1;
        layer_1_weights[539][8] = 0;
        layer_1_weights[540][8] = -1;
        layer_1_weights[541][8] = 2;
        layer_1_weights[542][8] = 1;
        layer_1_weights[543][8] = 2;
        layer_1_weights[544][8] = 1;
        layer_1_weights[545][8] = 1;
        layer_1_weights[546][8] = 1;
        layer_1_weights[547][8] = 2;
        layer_1_weights[548][8] = 1;
        layer_1_weights[549][8] = 1;
        layer_1_weights[550][8] = 1;
        layer_1_weights[551][8] = 0;
        layer_1_weights[552][8] = -1;
        layer_1_weights[553][8] = 0;
        layer_1_weights[554][8] = 2;
        layer_1_weights[555][8] = 1;
        layer_1_weights[556][8] = -1;
        layer_1_weights[557][8] = -1;
        layer_1_weights[558][8] = -5;
        layer_1_weights[559][8] = -3;
        layer_1_weights[560][8] = 0;
        layer_1_weights[561][8] = 2;
        layer_1_weights[562][8] = -2;
        layer_1_weights[563][8] = 1;
        layer_1_weights[564][8] = 2;
        layer_1_weights[565][8] = 1;
        layer_1_weights[566][8] = 0;
        layer_1_weights[567][8] = 1;
        layer_1_weights[568][8] = 0;
        layer_1_weights[569][8] = 0;
        layer_1_weights[570][8] = 1;
        layer_1_weights[571][8] = 3;
        layer_1_weights[572][8] = 2;
        layer_1_weights[573][8] = 1;
        layer_1_weights[574][8] = 2;
        layer_1_weights[575][8] = 2;
        layer_1_weights[576][8] = 2;
        layer_1_weights[577][8] = 1;
        layer_1_weights[578][8] = 1;
        layer_1_weights[579][8] = -1;
        layer_1_weights[580][8] = -1;
        layer_1_weights[581][8] = 2;
        layer_1_weights[582][8] = 0;
        layer_1_weights[583][8] = 1;
        layer_1_weights[584][8] = -5;
        layer_1_weights[585][8] = -3;
        layer_1_weights[586][8] = -4;
        layer_1_weights[587][8] = -2;
        layer_1_weights[588][8] = 0;
        layer_1_weights[589][8] = 1;
        layer_1_weights[590][8] = 1;
        layer_1_weights[591][8] = 2;
        layer_1_weights[592][8] = 1;
        layer_1_weights[593][8] = -2;
        layer_1_weights[594][8] = 0;
        layer_1_weights[595][8] = 1;
        layer_1_weights[596][8] = 0;
        layer_1_weights[597][8] = 1;
        layer_1_weights[598][8] = 1;
        layer_1_weights[599][8] = 1;
        layer_1_weights[600][8] = 1;
        layer_1_weights[601][8] = 1;
        layer_1_weights[602][8] = 2;
        layer_1_weights[603][8] = 1;
        layer_1_weights[604][8] = 1;
        layer_1_weights[605][8] = 1;
        layer_1_weights[606][8] = 1;
        layer_1_weights[607][8] = 0;
        layer_1_weights[608][8] = 0;
        layer_1_weights[609][8] = -2;
        layer_1_weights[610][8] = 0;
        layer_1_weights[611][8] = 0;
        layer_1_weights[612][8] = -3;
        layer_1_weights[613][8] = -1;
        layer_1_weights[614][8] = 2;
        layer_1_weights[615][8] = 1;
        layer_1_weights[616][8] = 0;
        layer_1_weights[617][8] = 1;
        layer_1_weights[618][8] = 1;
        layer_1_weights[619][8] = 0;
        layer_1_weights[620][8] = -1;
        layer_1_weights[621][8] = -2;
        layer_1_weights[622][8] = 0;
        layer_1_weights[623][8] = -2;
        layer_1_weights[624][8] = -1;
        layer_1_weights[625][8] = 0;
        layer_1_weights[626][8] = 0;
        layer_1_weights[627][8] = 3;
        layer_1_weights[628][8] = 1;
        layer_1_weights[629][8] = 2;
        layer_1_weights[630][8] = 1;
        layer_1_weights[631][8] = 1;
        layer_1_weights[632][8] = 1;
        layer_1_weights[633][8] = 1;
        layer_1_weights[634][8] = -1;
        layer_1_weights[635][8] = 1;
        layer_1_weights[636][8] = 0;
        layer_1_weights[637][8] = -2;
        layer_1_weights[638][8] = 1;
        layer_1_weights[639][8] = 2;
        layer_1_weights[640][8] = -2;
        layer_1_weights[641][8] = -1;
        layer_1_weights[642][8] = 4;
        layer_1_weights[643][8] = 1;
        layer_1_weights[644][8] = 0;
        layer_1_weights[645][8] = 0;
        layer_1_weights[646][8] = 3;
        layer_1_weights[647][8] = 5;
        layer_1_weights[648][8] = 4;
        layer_1_weights[649][8] = -2;
        layer_1_weights[650][8] = 1;
        layer_1_weights[651][8] = 0;
        layer_1_weights[652][8] = 2;
        layer_1_weights[653][8] = 0;
        layer_1_weights[654][8] = 0;
        layer_1_weights[655][8] = 0;
        layer_1_weights[656][8] = 1;
        layer_1_weights[657][8] = 1;
        layer_1_weights[658][8] = 1;
        layer_1_weights[659][8] = 1;
        layer_1_weights[660][8] = 0;
        layer_1_weights[661][8] = 2;
        layer_1_weights[662][8] = 1;
        layer_1_weights[663][8] = 2;
        layer_1_weights[664][8] = -2;
        layer_1_weights[665][8] = -1;
        layer_1_weights[666][8] = -1;
        layer_1_weights[667][8] = 1;
        layer_1_weights[668][8] = -1;
        layer_1_weights[669][8] = 1;
        layer_1_weights[670][8] = 2;
        layer_1_weights[671][8] = 0;
        layer_1_weights[672][8] = 1;
        layer_1_weights[673][8] = -1;
        layer_1_weights[674][8] = -2;
        layer_1_weights[675][8] = 2;
        layer_1_weights[676][8] = 0;
        layer_1_weights[677][8] = -1;
        layer_1_weights[678][8] = 1;
        layer_1_weights[679][8] = 0;
        layer_1_weights[680][8] = 1;
        layer_1_weights[681][8] = 0;
        layer_1_weights[682][8] = 2;
        layer_1_weights[683][8] = 1;
        layer_1_weights[684][8] = 2;
        layer_1_weights[685][8] = 2;
        layer_1_weights[686][8] = 3;
        layer_1_weights[687][8] = 1;
        layer_1_weights[688][8] = 1;
        layer_1_weights[689][8] = 0;
        layer_1_weights[690][8] = 2;
        layer_1_weights[691][8] = 0;
        layer_1_weights[692][8] = 1;
        layer_1_weights[693][8] = -3;
        layer_1_weights[694][8] = 2;
        layer_1_weights[695][8] = 1;
        layer_1_weights[696][8] = 1;
        layer_1_weights[697][8] = 2;
        layer_1_weights[698][8] = 0;
        layer_1_weights[699][8] = 0;
        layer_1_weights[700][8] = 0;
        layer_1_weights[701][8] = 1;
        layer_1_weights[702][8] = -1;
        layer_1_weights[703][8] = 1;
        layer_1_weights[704][8] = 0;
        layer_1_weights[705][8] = -1;
        layer_1_weights[706][8] = -2;
        layer_1_weights[707][8] = 1;
        layer_1_weights[708][8] = -3;
        layer_1_weights[709][8] = -1;
        layer_1_weights[710][8] = -1;
        layer_1_weights[711][8] = -1;
        layer_1_weights[712][8] = -2;
        layer_1_weights[713][8] = 0;
        layer_1_weights[714][8] = 0;
        layer_1_weights[715][8] = -1;
        layer_1_weights[716][8] = 0;
        layer_1_weights[717][8] = -2;
        layer_1_weights[718][8] = 0;
        layer_1_weights[719][8] = -3;
        layer_1_weights[720][8] = -1;
        layer_1_weights[721][8] = 0;
        layer_1_weights[722][8] = -2;
        layer_1_weights[723][8] = 1;
        layer_1_weights[724][8] = 2;
        layer_1_weights[725][8] = 0;
        layer_1_weights[726][8] = 0;
        layer_1_weights[727][8] = 0;
        layer_1_weights[728][8] = 0;
        layer_1_weights[729][8] = 1;
        layer_1_weights[730][8] = 0;
        layer_1_weights[731][8] = -3;
        layer_1_weights[732][8] = -1;
        layer_1_weights[733][8] = -2;
        layer_1_weights[734][8] = -3;
        layer_1_weights[735][8] = -7;
        layer_1_weights[736][8] = -3;
        layer_1_weights[737][8] = -5;
        layer_1_weights[738][8] = -4;
        layer_1_weights[739][8] = -3;
        layer_1_weights[740][8] = -3;
        layer_1_weights[741][8] = -2;
        layer_1_weights[742][8] = -3;
        layer_1_weights[743][8] = -5;
        layer_1_weights[744][8] = -2;
        layer_1_weights[745][8] = -3;
        layer_1_weights[746][8] = -3;
        layer_1_weights[747][8] = -2;
        layer_1_weights[748][8] = -3;
        layer_1_weights[749][8] = -5;
        layer_1_weights[750][8] = 0;
        layer_1_weights[751][8] = 0;
        layer_1_weights[752][8] = 0;
        layer_1_weights[753][8] = -1;
        layer_1_weights[754][8] = 0;
        layer_1_weights[755][8] = -1;
        layer_1_weights[756][8] = 0;
        layer_1_weights[757][8] = 0;
        layer_1_weights[758][8] = 0;
        layer_1_weights[759][8] = 0;
        layer_1_weights[760][8] = 0;
        layer_1_weights[761][8] = -1;
        layer_1_weights[762][8] = 0;
        layer_1_weights[763][8] = -2;
        layer_1_weights[764][8] = -3;
        layer_1_weights[765][8] = -5;
        layer_1_weights[766][8] = -4;
        layer_1_weights[767][8] = -3;
        layer_1_weights[768][8] = -2;
        layer_1_weights[769][8] = -3;
        layer_1_weights[770][8] = -8;
        layer_1_weights[771][8] = -3;
        layer_1_weights[772][8] = -2;
        layer_1_weights[773][8] = -4;
        layer_1_weights[774][8] = -2;
        layer_1_weights[775][8] = -2;
        layer_1_weights[776][8] = 1;
        layer_1_weights[777][8] = -1;
        layer_1_weights[778][8] = -2;
        layer_1_weights[779][8] = -1;
        layer_1_weights[780][8] = 0;
        layer_1_weights[781][8] = 1;
        layer_1_weights[782][8] = -1;
        layer_1_weights[783][8] = 0;
        layer_1_weights[0][9] = -1;
        layer_1_weights[1][9] = 0;
        layer_1_weights[2][9] = -1;
        layer_1_weights[3][9] = 0;
        layer_1_weights[4][9] = 1;
        layer_1_weights[5][9] = 0;
        layer_1_weights[6][9] = 0;
        layer_1_weights[7][9] = 0;
        layer_1_weights[8][9] = 1;
        layer_1_weights[9][9] = 0;
        layer_1_weights[10][9] = 0;
        layer_1_weights[11][9] = 0;
        layer_1_weights[12][9] = -1;
        layer_1_weights[13][9] = -1;
        layer_1_weights[14][9] = 2;
        layer_1_weights[15][9] = 1;
        layer_1_weights[16][9] = 0;
        layer_1_weights[17][9] = 1;
        layer_1_weights[18][9] = 1;
        layer_1_weights[19][9] = 0;
        layer_1_weights[20][9] = 0;
        layer_1_weights[21][9] = 0;
        layer_1_weights[22][9] = 0;
        layer_1_weights[23][9] = 1;
        layer_1_weights[24][9] = 0;
        layer_1_weights[25][9] = 1;
        layer_1_weights[26][9] = 0;
        layer_1_weights[27][9] = 0;
        layer_1_weights[28][9] = 0;
        layer_1_weights[29][9] = -1;
        layer_1_weights[30][9] = 0;
        layer_1_weights[31][9] = 0;
        layer_1_weights[32][9] = 0;
        layer_1_weights[33][9] = -3;
        layer_1_weights[34][9] = -2;
        layer_1_weights[35][9] = -4;
        layer_1_weights[36][9] = -4;
        layer_1_weights[37][9] = -4;
        layer_1_weights[38][9] = -6;
        layer_1_weights[39][9] = -6;
        layer_1_weights[40][9] = -5;
        layer_1_weights[41][9] = -6;
        layer_1_weights[42][9] = 2;
        layer_1_weights[43][9] = -4;
        layer_1_weights[44][9] = -3;
        layer_1_weights[45][9] = -4;
        layer_1_weights[46][9] = -6;
        layer_1_weights[47][9] = -5;
        layer_1_weights[48][9] = -4;
        layer_1_weights[49][9] = -4;
        layer_1_weights[50][9] = -2;
        layer_1_weights[51][9] = -2;
        layer_1_weights[52][9] = -1;
        layer_1_weights[53][9] = 0;
        layer_1_weights[54][9] = 0;
        layer_1_weights[55][9] = 1;
        layer_1_weights[56][9] = 0;
        layer_1_weights[57][9] = -1;
        layer_1_weights[58][9] = -2;
        layer_1_weights[59][9] = 0;
        layer_1_weights[60][9] = -3;
        layer_1_weights[61][9] = -2;
        layer_1_weights[62][9] = -4;
        layer_1_weights[63][9] = -6;
        layer_1_weights[64][9] = -7;
        layer_1_weights[65][9] = -5;
        layer_1_weights[66][9] = -7;
        layer_1_weights[67][9] = -7;
        layer_1_weights[68][9] = -4;
        layer_1_weights[69][9] = -1;
        layer_1_weights[70][9] = 0;
        layer_1_weights[71][9] = -1;
        layer_1_weights[72][9] = -3;
        layer_1_weights[73][9] = 0;
        layer_1_weights[74][9] = -1;
        layer_1_weights[75][9] = -3;
        layer_1_weights[76][9] = -1;
        layer_1_weights[77][9] = -2;
        layer_1_weights[78][9] = -1;
        layer_1_weights[79][9] = -2;
        layer_1_weights[80][9] = -4;
        layer_1_weights[81][9] = -2;
        layer_1_weights[82][9] = 1;
        layer_1_weights[83][9] = 0;
        layer_1_weights[84][9] = 1;
        layer_1_weights[85][9] = 0;
        layer_1_weights[86][9] = 2;
        layer_1_weights[87][9] = -2;
        layer_1_weights[88][9] = 1;
        layer_1_weights[89][9] = -3;
        layer_1_weights[90][9] = -5;
        layer_1_weights[91][9] = -1;
        layer_1_weights[92][9] = -4;
        layer_1_weights[93][9] = -5;
        layer_1_weights[94][9] = -4;
        layer_1_weights[95][9] = -2;
        layer_1_weights[96][9] = 0;
        layer_1_weights[97][9] = -2;
        layer_1_weights[98][9] = -1;
        layer_1_weights[99][9] = 1;
        layer_1_weights[100][9] = 1;
        layer_1_weights[101][9] = 0;
        layer_1_weights[102][9] = 1;
        layer_1_weights[103][9] = 0;
        layer_1_weights[104][9] = 0;
        layer_1_weights[105][9] = 1;
        layer_1_weights[106][9] = 2;
        layer_1_weights[107][9] = -1;
        layer_1_weights[108][9] = -1;
        layer_1_weights[109][9] = -3;
        layer_1_weights[110][9] = -3;
        layer_1_weights[111][9] = -1;
        layer_1_weights[112][9] = 0;
        layer_1_weights[113][9] = 2;
        layer_1_weights[114][9] = 2;
        layer_1_weights[115][9] = 0;
        layer_1_weights[116][9] = 0;
        layer_1_weights[117][9] = 1;
        layer_1_weights[118][9] = 1;
        layer_1_weights[119][9] = 1;
        layer_1_weights[120][9] = -3;
        layer_1_weights[121][9] = -1;
        layer_1_weights[122][9] = 0;
        layer_1_weights[123][9] = 1;
        layer_1_weights[124][9] = 1;
        layer_1_weights[125][9] = 1;
        layer_1_weights[126][9] = 2;
        layer_1_weights[127][9] = 2;
        layer_1_weights[128][9] = 0;
        layer_1_weights[129][9] = 0;
        layer_1_weights[130][9] = 0;
        layer_1_weights[131][9] = 1;
        layer_1_weights[132][9] = 0;
        layer_1_weights[133][9] = 1;
        layer_1_weights[134][9] = 0;
        layer_1_weights[135][9] = -1;
        layer_1_weights[136][9] = 2;
        layer_1_weights[137][9] = 1;
        layer_1_weights[138][9] = 2;
        layer_1_weights[139][9] = 0;
        layer_1_weights[140][9] = 0;
        layer_1_weights[141][9] = 1;
        layer_1_weights[142][9] = -3;
        layer_1_weights[143][9] = 6;
        layer_1_weights[144][9] = 2;
        layer_1_weights[145][9] = 3;
        layer_1_weights[146][9] = 2;
        layer_1_weights[147][9] = 0;
        layer_1_weights[148][9] = 0;
        layer_1_weights[149][9] = 0;
        layer_1_weights[150][9] = 0;
        layer_1_weights[151][9] = 2;
        layer_1_weights[152][9] = 0;
        layer_1_weights[153][9] = -2;
        layer_1_weights[154][9] = 2;
        layer_1_weights[155][9] = 1;
        layer_1_weights[156][9] = 1;
        layer_1_weights[157][9] = 0;
        layer_1_weights[158][9] = 0;
        layer_1_weights[159][9] = -2;
        layer_1_weights[160][9] = 2;
        layer_1_weights[161][9] = 0;
        layer_1_weights[162][9] = 0;
        layer_1_weights[163][9] = -1;
        layer_1_weights[164][9] = 2;
        layer_1_weights[165][9] = 4;
        layer_1_weights[166][9] = -1;
        layer_1_weights[167][9] = 1;
        layer_1_weights[168][9] = 0;
        layer_1_weights[169][9] = 1;
        layer_1_weights[170][9] = 1;
        layer_1_weights[171][9] = 3;
        layer_1_weights[172][9] = 1;
        layer_1_weights[173][9] = 0;
        layer_1_weights[174][9] = 1;
        layer_1_weights[175][9] = -1;
        layer_1_weights[176][9] = 3;
        layer_1_weights[177][9] = 2;
        layer_1_weights[178][9] = 0;
        layer_1_weights[179][9] = 0;
        layer_1_weights[180][9] = 1;
        layer_1_weights[181][9] = 0;
        layer_1_weights[182][9] = -1;
        layer_1_weights[183][9] = 0;
        layer_1_weights[184][9] = 0;
        layer_1_weights[185][9] = 0;
        layer_1_weights[186][9] = 1;
        layer_1_weights[187][9] = 1;
        layer_1_weights[188][9] = 2;
        layer_1_weights[189][9] = 0;
        layer_1_weights[190][9] = 0;
        layer_1_weights[191][9] = 0;
        layer_1_weights[192][9] = 4;
        layer_1_weights[193][9] = 0;
        layer_1_weights[194][9] = 1;
        layer_1_weights[195][9] = -1;
        layer_1_weights[196][9] = 0;
        layer_1_weights[197][9] = 2;
        layer_1_weights[198][9] = 0;
        layer_1_weights[199][9] = 4;
        layer_1_weights[200][9] = 5;
        layer_1_weights[201][9] = 2;
        layer_1_weights[202][9] = 0;
        layer_1_weights[203][9] = 1;
        layer_1_weights[204][9] = 2;
        layer_1_weights[205][9] = -1;
        layer_1_weights[206][9] = -2;
        layer_1_weights[207][9] = 0;
        layer_1_weights[208][9] = -1;
        layer_1_weights[209][9] = 0;
        layer_1_weights[210][9] = 0;
        layer_1_weights[211][9] = 0;
        layer_1_weights[212][9] = 1;
        layer_1_weights[213][9] = 0;
        layer_1_weights[214][9] = 0;
        layer_1_weights[215][9] = 1;
        layer_1_weights[216][9] = 2;
        layer_1_weights[217][9] = 2;
        layer_1_weights[218][9] = 0;
        layer_1_weights[219][9] = 0;
        layer_1_weights[220][9] = 0;
        layer_1_weights[221][9] = 1;
        layer_1_weights[222][9] = 5;
        layer_1_weights[223][9] = -1;
        layer_1_weights[224][9] = -3;
        layer_1_weights[225][9] = -4;
        layer_1_weights[226][9] = -1;
        layer_1_weights[227][9] = 0;
        layer_1_weights[228][9] = 3;
        layer_1_weights[229][9] = 3;
        layer_1_weights[230][9] = 1;
        layer_1_weights[231][9] = 2;
        layer_1_weights[232][9] = 2;
        layer_1_weights[233][9] = 2;
        layer_1_weights[234][9] = -1;
        layer_1_weights[235][9] = -1;
        layer_1_weights[236][9] = -1;
        layer_1_weights[237][9] = 0;
        layer_1_weights[238][9] = -1;
        layer_1_weights[239][9] = -1;
        layer_1_weights[240][9] = 0;
        layer_1_weights[241][9] = -2;
        layer_1_weights[242][9] = -1;
        layer_1_weights[243][9] = 1;
        layer_1_weights[244][9] = 1;
        layer_1_weights[245][9] = 0;
        layer_1_weights[246][9] = 2;
        layer_1_weights[247][9] = 1;
        layer_1_weights[248][9] = 0;
        layer_1_weights[249][9] = 3;
        layer_1_weights[250][9] = 2;
        layer_1_weights[251][9] = 2;
        layer_1_weights[252][9] = -3;
        layer_1_weights[253][9] = -2;
        layer_1_weights[254][9] = 2;
        layer_1_weights[255][9] = -1;
        layer_1_weights[256][9] = 1;
        layer_1_weights[257][9] = 2;
        layer_1_weights[258][9] = 1;
        layer_1_weights[259][9] = 1;
        layer_1_weights[260][9] = 0;
        layer_1_weights[261][9] = -1;
        layer_1_weights[262][9] = -2;
        layer_1_weights[263][9] = -1;
        layer_1_weights[264][9] = -1;
        layer_1_weights[265][9] = -1;
        layer_1_weights[266][9] = -1;
        layer_1_weights[267][9] = -1;
        layer_1_weights[268][9] = -1;
        layer_1_weights[269][9] = -1;
        layer_1_weights[270][9] = -1;
        layer_1_weights[271][9] = 0;
        layer_1_weights[272][9] = -1;
        layer_1_weights[273][9] = 0;
        layer_1_weights[274][9] = 0;
        layer_1_weights[275][9] = 1;
        layer_1_weights[276][9] = -1;
        layer_1_weights[277][9] = 5;
        layer_1_weights[278][9] = 4;
        layer_1_weights[279][9] = -2;
        layer_1_weights[280][9] = -2;
        layer_1_weights[281][9] = -2;
        layer_1_weights[282][9] = -2;
        layer_1_weights[283][9] = 0;
        layer_1_weights[284][9] = 3;
        layer_1_weights[285][9] = 0;
        layer_1_weights[286][9] = 0;
        layer_1_weights[287][9] = -2;
        layer_1_weights[288][9] = 1;
        layer_1_weights[289][9] = 0;
        layer_1_weights[290][9] = 1;
        layer_1_weights[291][9] = 0;
        layer_1_weights[292][9] = 0;
        layer_1_weights[293][9] = 0;
        layer_1_weights[294][9] = -1;
        layer_1_weights[295][9] = 0;
        layer_1_weights[296][9] = -2;
        layer_1_weights[297][9] = -2;
        layer_1_weights[298][9] = 0;
        layer_1_weights[299][9] = 0;
        layer_1_weights[300][9] = 1;
        layer_1_weights[301][9] = -1;
        layer_1_weights[302][9] = 0;
        layer_1_weights[303][9] = 0;
        layer_1_weights[304][9] = 0;
        layer_1_weights[305][9] = 2;
        layer_1_weights[306][9] = 0;
        layer_1_weights[307][9] = 1;
        layer_1_weights[308][9] = -2;
        layer_1_weights[309][9] = -4;
        layer_1_weights[310][9] = 1;
        layer_1_weights[311][9] = 2;
        layer_1_weights[312][9] = 2;
        layer_1_weights[313][9] = 0;
        layer_1_weights[314][9] = 1;
        layer_1_weights[315][9] = 0;
        layer_1_weights[316][9] = 2;
        layer_1_weights[317][9] = 1;
        layer_1_weights[318][9] = 1;
        layer_1_weights[319][9] = 1;
        layer_1_weights[320][9] = 2;
        layer_1_weights[321][9] = -1;
        layer_1_weights[322][9] = 0;
        layer_1_weights[323][9] = 1;
        layer_1_weights[324][9] = 0;
        layer_1_weights[325][9] = 0;
        layer_1_weights[326][9] = 0;
        layer_1_weights[327][9] = 0;
        layer_1_weights[328][9] = 0;
        layer_1_weights[329][9] = -2;
        layer_1_weights[330][9] = -2;
        layer_1_weights[331][9] = -2;
        layer_1_weights[332][9] = -2;
        layer_1_weights[333][9] = 1;
        layer_1_weights[334][9] = 2;
        layer_1_weights[335][9] = 2;
        layer_1_weights[336][9] = -1;
        layer_1_weights[337][9] = -4;
        layer_1_weights[338][9] = -3;
        layer_1_weights[339][9] = 0;
        layer_1_weights[340][9] = 0;
        layer_1_weights[341][9] = 1;
        layer_1_weights[342][9] = 1;
        layer_1_weights[343][9] = 1;
        layer_1_weights[344][9] = 2;
        layer_1_weights[345][9] = 1;
        layer_1_weights[346][9] = 3;
        layer_1_weights[347][9] = 2;
        layer_1_weights[348][9] = 2;
        layer_1_weights[349][9] = 1;
        layer_1_weights[350][9] = 1;
        layer_1_weights[351][9] = 2;
        layer_1_weights[352][9] = 2;
        layer_1_weights[353][9] = 3;
        layer_1_weights[354][9] = -1;
        layer_1_weights[355][9] = 2;
        layer_1_weights[356][9] = 0;
        layer_1_weights[357][9] = 0;
        layer_1_weights[358][9] = 0;
        layer_1_weights[359][9] = -2;
        layer_1_weights[360][9] = -3;
        layer_1_weights[361][9] = -1;
        layer_1_weights[362][9] = 2;
        layer_1_weights[363][9] = 3;
        layer_1_weights[364][9] = 0;
        layer_1_weights[365][9] = -2;
        layer_1_weights[366][9] = 0;
        layer_1_weights[367][9] = 2;
        layer_1_weights[368][9] = -1;
        layer_1_weights[369][9] = 0;
        layer_1_weights[370][9] = 1;
        layer_1_weights[371][9] = 1;
        layer_1_weights[372][9] = 3;
        layer_1_weights[373][9] = 2;
        layer_1_weights[374][9] = 2;
        layer_1_weights[375][9] = 2;
        layer_1_weights[376][9] = 2;
        layer_1_weights[377][9] = 2;
        layer_1_weights[378][9] = 4;
        layer_1_weights[379][9] = 2;
        layer_1_weights[380][9] = 4;
        layer_1_weights[381][9] = 3;
        layer_1_weights[382][9] = 1;
        layer_1_weights[383][9] = 2;
        layer_1_weights[384][9] = 1;
        layer_1_weights[385][9] = 0;
        layer_1_weights[386][9] = 0;
        layer_1_weights[387][9] = 0;
        layer_1_weights[388][9] = -3;
        layer_1_weights[389][9] = -1;
        layer_1_weights[390][9] = -1;
        layer_1_weights[391][9] = 2;
        layer_1_weights[392][9] = -1;
        layer_1_weights[393][9] = 1;
        layer_1_weights[394][9] = -3;
        layer_1_weights[395][9] = 3;
        layer_1_weights[396][9] = 1;
        layer_1_weights[397][9] = 1;
        layer_1_weights[398][9] = 0;
        layer_1_weights[399][9] = 1;
        layer_1_weights[400][9] = 2;
        layer_1_weights[401][9] = 1;
        layer_1_weights[402][9] = -1;
        layer_1_weights[403][9] = -1;
        layer_1_weights[404][9] = 1;
        layer_1_weights[405][9] = 1;
        layer_1_weights[406][9] = 4;
        layer_1_weights[407][9] = 4;
        layer_1_weights[408][9] = 5;
        layer_1_weights[409][9] = 2;
        layer_1_weights[410][9] = 1;
        layer_1_weights[411][9] = 1;
        layer_1_weights[412][9] = 0;
        layer_1_weights[413][9] = -1;
        layer_1_weights[414][9] = -2;
        layer_1_weights[415][9] = -1;
        layer_1_weights[416][9] = 0;
        layer_1_weights[417][9] = 0;
        layer_1_weights[418][9] = 1;
        layer_1_weights[419][9] = -1;
        layer_1_weights[420][9] = -2;
        layer_1_weights[421][9] = 2;
        layer_1_weights[422][9] = 4;
        layer_1_weights[423][9] = 7;
        layer_1_weights[424][9] = 0;
        layer_1_weights[425][9] = 0;
        layer_1_weights[426][9] = 0;
        layer_1_weights[427][9] = -1;
        layer_1_weights[428][9] = 0;
        layer_1_weights[429][9] = 0;
        layer_1_weights[430][9] = -1;
        layer_1_weights[431][9] = -1;
        layer_1_weights[432][9] = 1;
        layer_1_weights[433][9] = 1;
        layer_1_weights[434][9] = 4;
        layer_1_weights[435][9] = 4;
        layer_1_weights[436][9] = 3;
        layer_1_weights[437][9] = 2;
        layer_1_weights[438][9] = 0;
        layer_1_weights[439][9] = 0;
        layer_1_weights[440][9] = 0;
        layer_1_weights[441][9] = 1;
        layer_1_weights[442][9] = -1;
        layer_1_weights[443][9] = 1;
        layer_1_weights[444][9] = 0;
        layer_1_weights[445][9] = -1;
        layer_1_weights[446][9] = 3;
        layer_1_weights[447][9] = -1;
        layer_1_weights[448][9] = -2;
        layer_1_weights[449][9] = 3;
        layer_1_weights[450][9] = 0;
        layer_1_weights[451][9] = 4;
        layer_1_weights[452][9] = 0;
        layer_1_weights[453][9] = -2;
        layer_1_weights[454][9] = 0;
        layer_1_weights[455][9] = -2;
        layer_1_weights[456][9] = -2;
        layer_1_weights[457][9] = -1;
        layer_1_weights[458][9] = -3;
        layer_1_weights[459][9] = -2;
        layer_1_weights[460][9] = 0;
        layer_1_weights[461][9] = 4;
        layer_1_weights[462][9] = 4;
        layer_1_weights[463][9] = 3;
        layer_1_weights[464][9] = 2;
        layer_1_weights[465][9] = 3;
        layer_1_weights[466][9] = 2;
        layer_1_weights[467][9] = 0;
        layer_1_weights[468][9] = -1;
        layer_1_weights[469][9] = 0;
        layer_1_weights[470][9] = 0;
        layer_1_weights[471][9] = -1;
        layer_1_weights[472][9] = -1;
        layer_1_weights[473][9] = -2;
        layer_1_weights[474][9] = 1;
        layer_1_weights[475][9] = -3;
        layer_1_weights[476][9] = 0;
        layer_1_weights[477][9] = 3;
        layer_1_weights[478][9] = 1;
        layer_1_weights[479][9] = 2;
        layer_1_weights[480][9] = -2;
        layer_1_weights[481][9] = -2;
        layer_1_weights[482][9] = 0;
        layer_1_weights[483][9] = -1;
        layer_1_weights[484][9] = -3;
        layer_1_weights[485][9] = -4;
        layer_1_weights[486][9] = -5;
        layer_1_weights[487][9] = -2;
        layer_1_weights[488][9] = 0;
        layer_1_weights[489][9] = 2;
        layer_1_weights[490][9] = 3;
        layer_1_weights[491][9] = 3;
        layer_1_weights[492][9] = 2;
        layer_1_weights[493][9] = 1;
        layer_1_weights[494][9] = 1;
        layer_1_weights[495][9] = 0;
        layer_1_weights[496][9] = -2;
        layer_1_weights[497][9] = 0;
        layer_1_weights[498][9] = 0;
        layer_1_weights[499][9] = 1;
        layer_1_weights[500][9] = 0;
        layer_1_weights[501][9] = -4;
        layer_1_weights[502][9] = 0;
        layer_1_weights[503][9] = -3;
        layer_1_weights[504][9] = -2;
        layer_1_weights[505][9] = 0;
        layer_1_weights[506][9] = 1;
        layer_1_weights[507][9] = 3;
        layer_1_weights[508][9] = -2;
        layer_1_weights[509][9] = -1;
        layer_1_weights[510][9] = -1;
        layer_1_weights[511][9] = -2;
        layer_1_weights[512][9] = -3;
        layer_1_weights[513][9] = -3;
        layer_1_weights[514][9] = -4;
        layer_1_weights[515][9] = -2;
        layer_1_weights[516][9] = -2;
        layer_1_weights[517][9] = 2;
        layer_1_weights[518][9] = 3;
        layer_1_weights[519][9] = 3;
        layer_1_weights[520][9] = 2;
        layer_1_weights[521][9] = 0;
        layer_1_weights[522][9] = 1;
        layer_1_weights[523][9] = 1;
        layer_1_weights[524][9] = 0;
        layer_1_weights[525][9] = 2;
        layer_1_weights[526][9] = -1;
        layer_1_weights[527][9] = -1;
        layer_1_weights[528][9] = -1;
        layer_1_weights[529][9] = -3;
        layer_1_weights[530][9] = -2;
        layer_1_weights[531][9] = 2;
        layer_1_weights[532][9] = 0;
        layer_1_weights[533][9] = -3;
        layer_1_weights[534][9] = -1;
        layer_1_weights[535][9] = 1;
        layer_1_weights[536][9] = -1;
        layer_1_weights[537][9] = 0;
        layer_1_weights[538][9] = -2;
        layer_1_weights[539][9] = -1;
        layer_1_weights[540][9] = -2;
        layer_1_weights[541][9] = -3;
        layer_1_weights[542][9] = -4;
        layer_1_weights[543][9] = -4;
        layer_1_weights[544][9] = -4;
        layer_1_weights[545][9] = 0;
        layer_1_weights[546][9] = 2;
        layer_1_weights[547][9] = 2;
        layer_1_weights[548][9] = 1;
        layer_1_weights[549][9] = 0;
        layer_1_weights[550][9] = 1;
        layer_1_weights[551][9] = 2;
        layer_1_weights[552][9] = 0;
        layer_1_weights[553][9] = 0;
        layer_1_weights[554][9] = -1;
        layer_1_weights[555][9] = -1;
        layer_1_weights[556][9] = -3;
        layer_1_weights[557][9] = 3;
        layer_1_weights[558][9] = -1;
        layer_1_weights[559][9] = 2;
        layer_1_weights[560][9] = 1;
        layer_1_weights[561][9] = 1;
        layer_1_weights[562][9] = -1;
        layer_1_weights[563][9] = 2;
        layer_1_weights[564][9] = 0;
        layer_1_weights[565][9] = 0;
        layer_1_weights[566][9] = -2;
        layer_1_weights[567][9] = -2;
        layer_1_weights[568][9] = -2;
        layer_1_weights[569][9] = -2;
        layer_1_weights[570][9] = -3;
        layer_1_weights[571][9] = -3;
        layer_1_weights[572][9] = -3;
        layer_1_weights[573][9] = 0;
        layer_1_weights[574][9] = 1;
        layer_1_weights[575][9] = 1;
        layer_1_weights[576][9] = 1;
        layer_1_weights[577][9] = 2;
        layer_1_weights[578][9] = 1;
        layer_1_weights[579][9] = 1;
        layer_1_weights[580][9] = 0;
        layer_1_weights[581][9] = 0;
        layer_1_weights[582][9] = -1;
        layer_1_weights[583][9] = 1;
        layer_1_weights[584][9] = -2;
        layer_1_weights[585][9] = 2;
        layer_1_weights[586][9] = -2;
        layer_1_weights[587][9] = 3;
        layer_1_weights[588][9] = 0;
        layer_1_weights[589][9] = 2;
        layer_1_weights[590][9] = 2;
        layer_1_weights[591][9] = 2;
        layer_1_weights[592][9] = 0;
        layer_1_weights[593][9] = -1;
        layer_1_weights[594][9] = -1;
        layer_1_weights[595][9] = -1;
        layer_1_weights[596][9] = -1;
        layer_1_weights[597][9] = -2;
        layer_1_weights[598][9] = -1;
        layer_1_weights[599][9] = -1;
        layer_1_weights[600][9] = -1;
        layer_1_weights[601][9] = 0;
        layer_1_weights[602][9] = 1;
        layer_1_weights[603][9] = 1;
        layer_1_weights[604][9] = 1;
        layer_1_weights[605][9] = 0;
        layer_1_weights[606][9] = 0;
        layer_1_weights[607][9] = 0;
        layer_1_weights[608][9] = 1;
        layer_1_weights[609][9] = 1;
        layer_1_weights[610][9] = 1;
        layer_1_weights[611][9] = 0;
        layer_1_weights[612][9] = -2;
        layer_1_weights[613][9] = 0;
        layer_1_weights[614][9] = -3;
        layer_1_weights[615][9] = 0;
        layer_1_weights[616][9] = 0;
        layer_1_weights[617][9] = 2;
        layer_1_weights[618][9] = 1;
        layer_1_weights[619][9] = 2;
        layer_1_weights[620][9] = 0;
        layer_1_weights[621][9] = -2;
        layer_1_weights[622][9] = -1;
        layer_1_weights[623][9] = -1;
        layer_1_weights[624][9] = 0;
        layer_1_weights[625][9] = -1;
        layer_1_weights[626][9] = 1;
        layer_1_weights[627][9] = 0;
        layer_1_weights[628][9] = -1;
        layer_1_weights[629][9] = -1;
        layer_1_weights[630][9] = 1;
        layer_1_weights[631][9] = 1;
        layer_1_weights[632][9] = 1;
        layer_1_weights[633][9] = 1;
        layer_1_weights[634][9] = 0;
        layer_1_weights[635][9] = 2;
        layer_1_weights[636][9] = 2;
        layer_1_weights[637][9] = 3;
        layer_1_weights[638][9] = 0;
        layer_1_weights[639][9] = 0;
        layer_1_weights[640][9] = 3;
        layer_1_weights[641][9] = 1;
        layer_1_weights[642][9] = 0;
        layer_1_weights[643][9] = 0;
        layer_1_weights[644][9] = 0;
        layer_1_weights[645][9] = 0;
        layer_1_weights[646][9] = 2;
        layer_1_weights[647][9] = 4;
        layer_1_weights[648][9] = 5;
        layer_1_weights[649][9] = -1;
        layer_1_weights[650][9] = 1;
        layer_1_weights[651][9] = 1;
        layer_1_weights[652][9] = -1;
        layer_1_weights[653][9] = 0;
        layer_1_weights[654][9] = 1;
        layer_1_weights[655][9] = 0;
        layer_1_weights[656][9] = 0;
        layer_1_weights[657][9] = 0;
        layer_1_weights[658][9] = 0;
        layer_1_weights[659][9] = 1;
        layer_1_weights[660][9] = 0;
        layer_1_weights[661][9] = 1;
        layer_1_weights[662][9] = 2;
        layer_1_weights[663][9] = 4;
        layer_1_weights[664][9] = 2;
        layer_1_weights[665][9] = 1;
        layer_1_weights[666][9] = 0;
        layer_1_weights[667][9] = 1;
        layer_1_weights[668][9] = 2;
        layer_1_weights[669][9] = 4;
        layer_1_weights[670][9] = 5;
        layer_1_weights[671][9] = -1;
        layer_1_weights[672][9] = 0;
        layer_1_weights[673][9] = 0;
        layer_1_weights[674][9] = -1;
        layer_1_weights[675][9] = 1;
        layer_1_weights[676][9] = 2;
        layer_1_weights[677][9] = 3;
        layer_1_weights[678][9] = 2;
        layer_1_weights[679][9] = 1;
        layer_1_weights[680][9] = 1;
        layer_1_weights[681][9] = 1;
        layer_1_weights[682][9] = 2;
        layer_1_weights[683][9] = 2;
        layer_1_weights[684][9] = 0;
        layer_1_weights[685][9] = 1;
        layer_1_weights[686][9] = 0;
        layer_1_weights[687][9] = 2;
        layer_1_weights[688][9] = 0;
        layer_1_weights[689][9] = 3;
        layer_1_weights[690][9] = -1;
        layer_1_weights[691][9] = 2;
        layer_1_weights[692][9] = 4;
        layer_1_weights[693][9] = 3;
        layer_1_weights[694][9] = 2;
        layer_1_weights[695][9] = 5;
        layer_1_weights[696][9] = -1;
        layer_1_weights[697][9] = 1;
        layer_1_weights[698][9] = -2;
        layer_1_weights[699][9] = 1;
        layer_1_weights[700][9] = 0;
        layer_1_weights[701][9] = 1;
        layer_1_weights[702][9] = 3;
        layer_1_weights[703][9] = -4;
        layer_1_weights[704][9] = 2;
        layer_1_weights[705][9] = 6;
        layer_1_weights[706][9] = 4;
        layer_1_weights[707][9] = 6;
        layer_1_weights[708][9] = 5;
        layer_1_weights[709][9] = 6;
        layer_1_weights[710][9] = 3;
        layer_1_weights[711][9] = 3;
        layer_1_weights[712][9] = 3;
        layer_1_weights[713][9] = 3;
        layer_1_weights[714][9] = 3;
        layer_1_weights[715][9] = 3;
        layer_1_weights[716][9] = 3;
        layer_1_weights[717][9] = 2;
        layer_1_weights[718][9] = 3;
        layer_1_weights[719][9] = 5;
        layer_1_weights[720][9] = 3;
        layer_1_weights[721][9] = 5;
        layer_1_weights[722][9] = 4;
        layer_1_weights[723][9] = 5;
        layer_1_weights[724][9] = -1;
        layer_1_weights[725][9] = 1;
        layer_1_weights[726][9] = -2;
        layer_1_weights[727][9] = -1;
        layer_1_weights[728][9] = 0;
        layer_1_weights[729][9] = 0;
        layer_1_weights[730][9] = 0;
        layer_1_weights[731][9] = -1;
        layer_1_weights[732][9] = 3;
        layer_1_weights[733][9] = 4;
        layer_1_weights[734][9] = 4;
        layer_1_weights[735][9] = 3;
        layer_1_weights[736][9] = 2;
        layer_1_weights[737][9] = 3;
        layer_1_weights[738][9] = 2;
        layer_1_weights[739][9] = 2;
        layer_1_weights[740][9] = 0;
        layer_1_weights[741][9] = 0;
        layer_1_weights[742][9] = 1;
        layer_1_weights[743][9] = 0;
        layer_1_weights[744][9] = 1;
        layer_1_weights[745][9] = 2;
        layer_1_weights[746][9] = 2;
        layer_1_weights[747][9] = -4;
        layer_1_weights[748][9] = -1;
        layer_1_weights[749][9] = 1;
        layer_1_weights[750][9] = -1;
        layer_1_weights[751][9] = -1;
        layer_1_weights[752][9] = 0;
        layer_1_weights[753][9] = -2;
        layer_1_weights[754][9] = 0;
        layer_1_weights[755][9] = 0;
        layer_1_weights[756][9] = 0;
        layer_1_weights[757][9] = 0;
        layer_1_weights[758][9] = 0;
        layer_1_weights[759][9] = 0;
        layer_1_weights[760][9] = -1;
        layer_1_weights[761][9] = -4;
        layer_1_weights[762][9] = 2;
        layer_1_weights[763][9] = 1;
        layer_1_weights[764][9] = 0;
        layer_1_weights[765][9] = -1;
        layer_1_weights[766][9] = -3;
        layer_1_weights[767][9] = -1;
        layer_1_weights[768][9] = -2;
        layer_1_weights[769][9] = -4;
        layer_1_weights[770][9] = -6;
        layer_1_weights[771][9] = 0;
        layer_1_weights[772][9] = 0;
        layer_1_weights[773][9] = -5;
        layer_1_weights[774][9] = -1;
        layer_1_weights[775][9] = -3;
        layer_1_weights[776][9] = 0;
        layer_1_weights[777][9] = -2;
        layer_1_weights[778][9] = -1;
        layer_1_weights[779][9] = -2;
        layer_1_weights[780][9] = 0;
        layer_1_weights[781][9] = -1;
        layer_1_weights[782][9] = 0;
        layer_1_weights[783][9] = 0;
        layer_1_weights[0][10] = 0;
        layer_1_weights[1][10] = 1;
        layer_1_weights[2][10] = 0;
        layer_1_weights[3][10] = 0;
        layer_1_weights[4][10] = 0;
        layer_1_weights[5][10] = -1;
        layer_1_weights[6][10] = 0;
        layer_1_weights[7][10] = 0;
        layer_1_weights[8][10] = 1;
        layer_1_weights[9][10] = 0;
        layer_1_weights[10][10] = 0;
        layer_1_weights[11][10] = 0;
        layer_1_weights[12][10] = -1;
        layer_1_weights[13][10] = -1;
        layer_1_weights[14][10] = -1;
        layer_1_weights[15][10] = 1;
        layer_1_weights[16][10] = 0;
        layer_1_weights[17][10] = 0;
        layer_1_weights[18][10] = 0;
        layer_1_weights[19][10] = 0;
        layer_1_weights[20][10] = 0;
        layer_1_weights[21][10] = 0;
        layer_1_weights[22][10] = 1;
        layer_1_weights[23][10] = 0;
        layer_1_weights[24][10] = 0;
        layer_1_weights[25][10] = 1;
        layer_1_weights[26][10] = 0;
        layer_1_weights[27][10] = 0;
        layer_1_weights[28][10] = 0;
        layer_1_weights[29][10] = 0;
        layer_1_weights[30][10] = 0;
        layer_1_weights[31][10] = 0;
        layer_1_weights[32][10] = -1;
        layer_1_weights[33][10] = -3;
        layer_1_weights[34][10] = -2;
        layer_1_weights[35][10] = -2;
        layer_1_weights[36][10] = -3;
        layer_1_weights[37][10] = -2;
        layer_1_weights[38][10] = -4;
        layer_1_weights[39][10] = 1;
        layer_1_weights[40][10] = 0;
        layer_1_weights[41][10] = 1;
        layer_1_weights[42][10] = 2;
        layer_1_weights[43][10] = -1;
        layer_1_weights[44][10] = -1;
        layer_1_weights[45][10] = 1;
        layer_1_weights[46][10] = -6;
        layer_1_weights[47][10] = -5;
        layer_1_weights[48][10] = -3;
        layer_1_weights[49][10] = -3;
        layer_1_weights[50][10] = -3;
        layer_1_weights[51][10] = -2;
        layer_1_weights[52][10] = -1;
        layer_1_weights[53][10] = -1;
        layer_1_weights[54][10] = 0;
        layer_1_weights[55][10] = 0;
        layer_1_weights[56][10] = 0;
        layer_1_weights[57][10] = 0;
        layer_1_weights[58][10] = -1;
        layer_1_weights[59][10] = 0;
        layer_1_weights[60][10] = -2;
        layer_1_weights[61][10] = -1;
        layer_1_weights[62][10] = 0;
        layer_1_weights[63][10] = -3;
        layer_1_weights[64][10] = -5;
        layer_1_weights[65][10] = -6;
        layer_1_weights[66][10] = -7;
        layer_1_weights[67][10] = -3;
        layer_1_weights[68][10] = -5;
        layer_1_weights[69][10] = 0;
        layer_1_weights[70][10] = -2;
        layer_1_weights[71][10] = -2;
        layer_1_weights[72][10] = -3;
        layer_1_weights[73][10] = -2;
        layer_1_weights[74][10] = -5;
        layer_1_weights[75][10] = -3;
        layer_1_weights[76][10] = -6;
        layer_1_weights[77][10] = -5;
        layer_1_weights[78][10] = -2;
        layer_1_weights[79][10] = -6;
        layer_1_weights[80][10] = -4;
        layer_1_weights[81][10] = -3;
        layer_1_weights[82][10] = 0;
        layer_1_weights[83][10] = 1;
        layer_1_weights[84][10] = 0;
        layer_1_weights[85][10] = 0;
        layer_1_weights[86][10] = -1;
        layer_1_weights[87][10] = -1;
        layer_1_weights[88][10] = -3;
        layer_1_weights[89][10] = -4;
        layer_1_weights[90][10] = -6;
        layer_1_weights[91][10] = -5;
        layer_1_weights[92][10] = -4;
        layer_1_weights[93][10] = -4;
        layer_1_weights[94][10] = -3;
        layer_1_weights[95][10] = -4;
        layer_1_weights[96][10] = -4;
        layer_1_weights[97][10] = -5;
        layer_1_weights[98][10] = -1;
        layer_1_weights[99][10] = -1;
        layer_1_weights[100][10] = 1;
        layer_1_weights[101][10] = 2;
        layer_1_weights[102][10] = 0;
        layer_1_weights[103][10] = -2;
        layer_1_weights[104][10] = 1;
        layer_1_weights[105][10] = -2;
        layer_1_weights[106][10] = -2;
        layer_1_weights[107][10] = -2;
        layer_1_weights[108][10] = -2;
        layer_1_weights[109][10] = -1;
        layer_1_weights[110][10] = 0;
        layer_1_weights[111][10] = 0;
        layer_1_weights[112][10] = 1;
        layer_1_weights[113][10] = 0;
        layer_1_weights[114][10] = 0;
        layer_1_weights[115][10] = 1;
        layer_1_weights[116][10] = -2;
        layer_1_weights[117][10] = -2;
        layer_1_weights[118][10] = 0;
        layer_1_weights[119][10] = 0;
        layer_1_weights[120][10] = -1;
        layer_1_weights[121][10] = -3;
        layer_1_weights[122][10] = -3;
        layer_1_weights[123][10] = -1;
        layer_1_weights[124][10] = -1;
        layer_1_weights[125][10] = 0;
        layer_1_weights[126][10] = -1;
        layer_1_weights[127][10] = 1;
        layer_1_weights[128][10] = -2;
        layer_1_weights[129][10] = -1;
        layer_1_weights[130][10] = 1;
        layer_1_weights[131][10] = -1;
        layer_1_weights[132][10] = 1;
        layer_1_weights[133][10] = -1;
        layer_1_weights[134][10] = 2;
        layer_1_weights[135][10] = 2;
        layer_1_weights[136][10] = 3;
        layer_1_weights[137][10] = 2;
        layer_1_weights[138][10] = 3;
        layer_1_weights[139][10] = 1;
        layer_1_weights[140][10] = 0;
        layer_1_weights[141][10] = -1;
        layer_1_weights[142][10] = -4;
        layer_1_weights[143][10] = 0;
        layer_1_weights[144][10] = -2;
        layer_1_weights[145][10] = 1;
        layer_1_weights[146][10] = 0;
        layer_1_weights[147][10] = 0;
        layer_1_weights[148][10] = 0;
        layer_1_weights[149][10] = 0;
        layer_1_weights[150][10] = 0;
        layer_1_weights[151][10] = 0;
        layer_1_weights[152][10] = 0;
        layer_1_weights[153][10] = 0;
        layer_1_weights[154][10] = 1;
        layer_1_weights[155][10] = -1;
        layer_1_weights[156][10] = 0;
        layer_1_weights[157][10] = 0;
        layer_1_weights[158][10] = 0;
        layer_1_weights[159][10] = 0;
        layer_1_weights[160][10] = 1;
        layer_1_weights[161][10] = 0;
        layer_1_weights[162][10] = 0;
        layer_1_weights[163][10] = -2;
        layer_1_weights[164][10] = -4;
        layer_1_weights[165][10] = 2;
        layer_1_weights[166][10] = -4;
        layer_1_weights[167][10] = -1;
        layer_1_weights[168][10] = 0;
        layer_1_weights[169][10] = -1;
        layer_1_weights[170][10] = 0;
        layer_1_weights[171][10] = 2;
        layer_1_weights[172][10] = -1;
        layer_1_weights[173][10] = 2;
        layer_1_weights[174][10] = 0;
        layer_1_weights[175][10] = 0;
        layer_1_weights[176][10] = -2;
        layer_1_weights[177][10] = 0;
        layer_1_weights[178][10] = 0;
        layer_1_weights[179][10] = 1;
        layer_1_weights[180][10] = 2;
        layer_1_weights[181][10] = 2;
        layer_1_weights[182][10] = -1;
        layer_1_weights[183][10] = 1;
        layer_1_weights[184][10] = 2;
        layer_1_weights[185][10] = 2;
        layer_1_weights[186][10] = 3;
        layer_1_weights[187][10] = 2;
        layer_1_weights[188][10] = 1;
        layer_1_weights[189][10] = 3;
        layer_1_weights[190][10] = 1;
        layer_1_weights[191][10] = 1;
        layer_1_weights[192][10] = -2;
        layer_1_weights[193][10] = -4;
        layer_1_weights[194][10] = -3;
        layer_1_weights[195][10] = -1;
        layer_1_weights[196][10] = 1;
        layer_1_weights[197][10] = -4;
        layer_1_weights[198][10] = 2;
        layer_1_weights[199][10] = 0;
        layer_1_weights[200][10] = -3;
        layer_1_weights[201][10] = 1;
        layer_1_weights[202][10] = 1;
        layer_1_weights[203][10] = -1;
        layer_1_weights[204][10] = 0;
        layer_1_weights[205][10] = 2;
        layer_1_weights[206][10] = 2;
        layer_1_weights[207][10] = 0;
        layer_1_weights[208][10] = 1;
        layer_1_weights[209][10] = 1;
        layer_1_weights[210][10] = 1;
        layer_1_weights[211][10] = 3;
        layer_1_weights[212][10] = 2;
        layer_1_weights[213][10] = 3;
        layer_1_weights[214][10] = 4;
        layer_1_weights[215][10] = 3;
        layer_1_weights[216][10] = 3;
        layer_1_weights[217][10] = 1;
        layer_1_weights[218][10] = 0;
        layer_1_weights[219][10] = 3;
        layer_1_weights[220][10] = 1;
        layer_1_weights[221][10] = -1;
        layer_1_weights[222][10] = -3;
        layer_1_weights[223][10] = -1;
        layer_1_weights[224][10] = 2;
        layer_1_weights[225][10] = -2;
        layer_1_weights[226][10] = 2;
        layer_1_weights[227][10] = 3;
        layer_1_weights[228][10] = 3;
        layer_1_weights[229][10] = -1;
        layer_1_weights[230][10] = 2;
        layer_1_weights[231][10] = -1;
        layer_1_weights[232][10] = 1;
        layer_1_weights[233][10] = 0;
        layer_1_weights[234][10] = 1;
        layer_1_weights[235][10] = 1;
        layer_1_weights[236][10] = 2;
        layer_1_weights[237][10] = 2;
        layer_1_weights[238][10] = 1;
        layer_1_weights[239][10] = 1;
        layer_1_weights[240][10] = 1;
        layer_1_weights[241][10] = 2;
        layer_1_weights[242][10] = 2;
        layer_1_weights[243][10] = 1;
        layer_1_weights[244][10] = 1;
        layer_1_weights[245][10] = 1;
        layer_1_weights[246][10] = 2;
        layer_1_weights[247][10] = 1;
        layer_1_weights[248][10] = 3;
        layer_1_weights[249][10] = -1;
        layer_1_weights[250][10] = -2;
        layer_1_weights[251][10] = -1;
        layer_1_weights[252][10] = 2;
        layer_1_weights[253][10] = 2;
        layer_1_weights[254][10] = 0;
        layer_1_weights[255][10] = 0;
        layer_1_weights[256][10] = 0;
        layer_1_weights[257][10] = 0;
        layer_1_weights[258][10] = 1;
        layer_1_weights[259][10] = 1;
        layer_1_weights[260][10] = 1;
        layer_1_weights[261][10] = 1;
        layer_1_weights[262][10] = 0;
        layer_1_weights[263][10] = 2;
        layer_1_weights[264][10] = 1;
        layer_1_weights[265][10] = 1;
        layer_1_weights[266][10] = 0;
        layer_1_weights[267][10] = 0;
        layer_1_weights[268][10] = 1;
        layer_1_weights[269][10] = 1;
        layer_1_weights[270][10] = 2;
        layer_1_weights[271][10] = 4;
        layer_1_weights[272][10] = 2;
        layer_1_weights[273][10] = 2;
        layer_1_weights[274][10] = 2;
        layer_1_weights[275][10] = 0;
        layer_1_weights[276][10] = 4;
        layer_1_weights[277][10] = -1;
        layer_1_weights[278][10] = -3;
        layer_1_weights[279][10] = 2;
        layer_1_weights[280][10] = 1;
        layer_1_weights[281][10] = 1;
        layer_1_weights[282][10] = 1;
        layer_1_weights[283][10] = 1;
        layer_1_weights[284][10] = 1;
        layer_1_weights[285][10] = -1;
        layer_1_weights[286][10] = 0;
        layer_1_weights[287][10] = 1;
        layer_1_weights[288][10] = 0;
        layer_1_weights[289][10] = 0;
        layer_1_weights[290][10] = 0;
        layer_1_weights[291][10] = 0;
        layer_1_weights[292][10] = -1;
        layer_1_weights[293][10] = 1;
        layer_1_weights[294][10] = -1;
        layer_1_weights[295][10] = -1;
        layer_1_weights[296][10] = -1;
        layer_1_weights[297][10] = 0;
        layer_1_weights[298][10] = 2;
        layer_1_weights[299][10] = 1;
        layer_1_weights[300][10] = 1;
        layer_1_weights[301][10] = 1;
        layer_1_weights[302][10] = 2;
        layer_1_weights[303][10] = 3;
        layer_1_weights[304][10] = 0;
        layer_1_weights[305][10] = -3;
        layer_1_weights[306][10] = -4;
        layer_1_weights[307][10] = 2;
        layer_1_weights[308][10] = 2;
        layer_1_weights[309][10] = 4;
        layer_1_weights[310][10] = 2;
        layer_1_weights[311][10] = 0;
        layer_1_weights[312][10] = -1;
        layer_1_weights[313][10] = 1;
        layer_1_weights[314][10] = 2;
        layer_1_weights[315][10] = 3;
        layer_1_weights[316][10] = 2;
        layer_1_weights[317][10] = 1;
        layer_1_weights[318][10] = 1;
        layer_1_weights[319][10] = 0;
        layer_1_weights[320][10] = 0;
        layer_1_weights[321][10] = -1;
        layer_1_weights[322][10] = 0;
        layer_1_weights[323][10] = -1;
        layer_1_weights[324][10] = 1;
        layer_1_weights[325][10] = 1;
        layer_1_weights[326][10] = 0;
        layer_1_weights[327][10] = 1;
        layer_1_weights[328][10] = 1;
        layer_1_weights[329][10] = 2;
        layer_1_weights[330][10] = 3;
        layer_1_weights[331][10] = 2;
        layer_1_weights[332][10] = 0;
        layer_1_weights[333][10] = -4;
        layer_1_weights[334][10] = -1;
        layer_1_weights[335][10] = 1;
        layer_1_weights[336][10] = 2;
        layer_1_weights[337][10] = 6;
        layer_1_weights[338][10] = 4;
        layer_1_weights[339][10] = 2;
        layer_1_weights[340][10] = 2;
        layer_1_weights[341][10] = 1;
        layer_1_weights[342][10] = 3;
        layer_1_weights[343][10] = 3;
        layer_1_weights[344][10] = 1;
        layer_1_weights[345][10] = 0;
        layer_1_weights[346][10] = 0;
        layer_1_weights[347][10] = 1;
        layer_1_weights[348][10] = -2;
        layer_1_weights[349][10] = 1;
        layer_1_weights[350][10] = -1;
        layer_1_weights[351][10] = 1;
        layer_1_weights[352][10] = 0;
        layer_1_weights[353][10] = 0;
        layer_1_weights[354][10] = 0;
        layer_1_weights[355][10] = 1;
        layer_1_weights[356][10] = 2;
        layer_1_weights[357][10] = 2;
        layer_1_weights[358][10] = 3;
        layer_1_weights[359][10] = 2;
        layer_1_weights[360][10] = 2;
        layer_1_weights[361][10] = -2;
        layer_1_weights[362][10] = -2;
        layer_1_weights[363][10] = 3;
        layer_1_weights[364][10] = 0;
        layer_1_weights[365][10] = 4;
        layer_1_weights[366][10] = 2;
        layer_1_weights[367][10] = 0;
        layer_1_weights[368][10] = 5;
        layer_1_weights[369][10] = 2;
        layer_1_weights[370][10] = 1;
        layer_1_weights[371][10] = 1;
        layer_1_weights[372][10] = 1;
        layer_1_weights[373][10] = -2;
        layer_1_weights[374][10] = 0;
        layer_1_weights[375][10] = -1;
        layer_1_weights[376][10] = -2;
        layer_1_weights[377][10] = -1;
        layer_1_weights[378][10] = 0;
        layer_1_weights[379][10] = 1;
        layer_1_weights[380][10] = 1;
        layer_1_weights[381][10] = -1;
        layer_1_weights[382][10] = 1;
        layer_1_weights[383][10] = 0;
        layer_1_weights[384][10] = 2;
        layer_1_weights[385][10] = 1;
        layer_1_weights[386][10] = 3;
        layer_1_weights[387][10] = 0;
        layer_1_weights[388][10] = -1;
        layer_1_weights[389][10] = 0;
        layer_1_weights[390][10] = -4;
        layer_1_weights[391][10] = -1;
        layer_1_weights[392][10] = -3;
        layer_1_weights[393][10] = 1;
        layer_1_weights[394][10] = 4;
        layer_1_weights[395][10] = -2;
        layer_1_weights[396][10] = 0;
        layer_1_weights[397][10] = 2;
        layer_1_weights[398][10] = 0;
        layer_1_weights[399][10] = 1;
        layer_1_weights[400][10] = 0;
        layer_1_weights[401][10] = 2;
        layer_1_weights[402][10] = 0;
        layer_1_weights[403][10] = 0;
        layer_1_weights[404][10] = 0;
        layer_1_weights[405][10] = 0;
        layer_1_weights[406][10] = 0;
        layer_1_weights[407][10] = 0;
        layer_1_weights[408][10] = 0;
        layer_1_weights[409][10] = 0;
        layer_1_weights[410][10] = 1;
        layer_1_weights[411][10] = 2;
        layer_1_weights[412][10] = 2;
        layer_1_weights[413][10] = 2;
        layer_1_weights[414][10] = 2;
        layer_1_weights[415][10] = 1;
        layer_1_weights[416][10] = 0;
        layer_1_weights[417][10] = 0;
        layer_1_weights[418][10] = -1;
        layer_1_weights[419][10] = 0;
        layer_1_weights[420][10] = -2;
        layer_1_weights[421][10] = 1;
        layer_1_weights[422][10] = -2;
        layer_1_weights[423][10] = -2;
        layer_1_weights[424][10] = 0;
        layer_1_weights[425][10] = 1;
        layer_1_weights[426][10] = 1;
        layer_1_weights[427][10] = 2;
        layer_1_weights[428][10] = 2;
        layer_1_weights[429][10] = 0;
        layer_1_weights[430][10] = 0;
        layer_1_weights[431][10] = 0;
        layer_1_weights[432][10] = 0;
        layer_1_weights[433][10] = 0;
        layer_1_weights[434][10] = -2;
        layer_1_weights[435][10] = 0;
        layer_1_weights[436][10] = -2;
        layer_1_weights[437][10] = -1;
        layer_1_weights[438][10] = 1;
        layer_1_weights[439][10] = 0;
        layer_1_weights[440][10] = 2;
        layer_1_weights[441][10] = 0;
        layer_1_weights[442][10] = 1;
        layer_1_weights[443][10] = 0;
        layer_1_weights[444][10] = -1;
        layer_1_weights[445][10] = -2;
        layer_1_weights[446][10] = -3;
        layer_1_weights[447][10] = -4;
        layer_1_weights[448][10] = 2;
        layer_1_weights[449][10] = 0;
        layer_1_weights[450][10] = 0;
        layer_1_weights[451][10] = -5;
        layer_1_weights[452][10] = 0;
        layer_1_weights[453][10] = 0;
        layer_1_weights[454][10] = 1;
        layer_1_weights[455][10] = 3;
        layer_1_weights[456][10] = 3;
        layer_1_weights[457][10] = 0;
        layer_1_weights[458][10] = 1;
        layer_1_weights[459][10] = 0;
        layer_1_weights[460][10] = 1;
        layer_1_weights[461][10] = 0;
        layer_1_weights[462][10] = -1;
        layer_1_weights[463][10] = 0;
        layer_1_weights[464][10] = 1;
        layer_1_weights[465][10] = 0;
        layer_1_weights[466][10] = -1;
        layer_1_weights[467][10] = 0;
        layer_1_weights[468][10] = 1;
        layer_1_weights[469][10] = -1;
        layer_1_weights[470][10] = 0;
        layer_1_weights[471][10] = -1;
        layer_1_weights[472][10] = 0;
        layer_1_weights[473][10] = -3;
        layer_1_weights[474][10] = -3;
        layer_1_weights[475][10] = -4;
        layer_1_weights[476][10] = 0;
        layer_1_weights[477][10] = -2;
        layer_1_weights[478][10] = 0;
        layer_1_weights[479][10] = -3;
        layer_1_weights[480][10] = 1;
        layer_1_weights[481][10] = 0;
        layer_1_weights[482][10] = 1;
        layer_1_weights[483][10] = 2;
        layer_1_weights[484][10] = 2;
        layer_1_weights[485][10] = 2;
        layer_1_weights[486][10] = 1;
        layer_1_weights[487][10] = 0;
        layer_1_weights[488][10] = 0;
        layer_1_weights[489][10] = -1;
        layer_1_weights[490][10] = 0;
        layer_1_weights[491][10] = 0;
        layer_1_weights[492][10] = 1;
        layer_1_weights[493][10] = 1;
        layer_1_weights[494][10] = 0;
        layer_1_weights[495][10] = 0;
        layer_1_weights[496][10] = 0;
        layer_1_weights[497][10] = 0;
        layer_1_weights[498][10] = 1;
        layer_1_weights[499][10] = 0;
        layer_1_weights[500][10] = 0;
        layer_1_weights[501][10] = -2;
        layer_1_weights[502][10] = -2;
        layer_1_weights[503][10] = 1;
        layer_1_weights[504][10] = 3;
        layer_1_weights[505][10] = 1;
        layer_1_weights[506][10] = 3;
        layer_1_weights[507][10] = -3;
        layer_1_weights[508][10] = -3;
        layer_1_weights[509][10] = -1;
        layer_1_weights[510][10] = -1;
        layer_1_weights[511][10] = -1;
        layer_1_weights[512][10] = 1;
        layer_1_weights[513][10] = 1;
        layer_1_weights[514][10] = 1;
        layer_1_weights[515][10] = -1;
        layer_1_weights[516][10] = -1;
        layer_1_weights[517][10] = 0;
        layer_1_weights[518][10] = 1;
        layer_1_weights[519][10] = 0;
        layer_1_weights[520][10] = 1;
        layer_1_weights[521][10] = 1;
        layer_1_weights[522][10] = -1;
        layer_1_weights[523][10] = -1;
        layer_1_weights[524][10] = 0;
        layer_1_weights[525][10] = 0;
        layer_1_weights[526][10] = -1;
        layer_1_weights[527][10] = -1;
        layer_1_weights[528][10] = -1;
        layer_1_weights[529][10] = -3;
        layer_1_weights[530][10] = -5;
        layer_1_weights[531][10] = -4;
        layer_1_weights[532][10] = 0;
        layer_1_weights[533][10] = 2;
        layer_1_weights[534][10] = 3;
        layer_1_weights[535][10] = -1;
        layer_1_weights[536][10] = 0;
        layer_1_weights[537][10] = -1;
        layer_1_weights[538][10] = 0;
        layer_1_weights[539][10] = -1;
        layer_1_weights[540][10] = -1;
        layer_1_weights[541][10] = -2;
        layer_1_weights[542][10] = -1;
        layer_1_weights[543][10] = -2;
        layer_1_weights[544][10] = -1;
        layer_1_weights[545][10] = -2;
        layer_1_weights[546][10] = 0;
        layer_1_weights[547][10] = 0;
        layer_1_weights[548][10] = 1;
        layer_1_weights[549][10] = 0;
        layer_1_weights[550][10] = 0;
        layer_1_weights[551][10] = 0;
        layer_1_weights[552][10] = 0;
        layer_1_weights[553][10] = 0;
        layer_1_weights[554][10] = 0;
        layer_1_weights[555][10] = -2;
        layer_1_weights[556][10] = -2;
        layer_1_weights[557][10] = -3;
        layer_1_weights[558][10] = -2;
        layer_1_weights[559][10] = -2;
        layer_1_weights[560][10] = 0;
        layer_1_weights[561][10] = 2;
        layer_1_weights[562][10] = -3;
        layer_1_weights[563][10] = -1;
        layer_1_weights[564][10] = 1;
        layer_1_weights[565][10] = 1;
        layer_1_weights[566][10] = -1;
        layer_1_weights[567][10] = -1;
        layer_1_weights[568][10] = -1;
        layer_1_weights[569][10] = -2;
        layer_1_weights[570][10] = -1;
        layer_1_weights[571][10] = -2;
        layer_1_weights[572][10] = -1;
        layer_1_weights[573][10] = -1;
        layer_1_weights[574][10] = 0;
        layer_1_weights[575][10] = -1;
        layer_1_weights[576][10] = -1;
        layer_1_weights[577][10] = 0;
        layer_1_weights[578][10] = -1;
        layer_1_weights[579][10] = -1;
        layer_1_weights[580][10] = -2;
        layer_1_weights[581][10] = 0;
        layer_1_weights[582][10] = -1;
        layer_1_weights[583][10] = -2;
        layer_1_weights[584][10] = 1;
        layer_1_weights[585][10] = 1;
        layer_1_weights[586][10] = -3;
        layer_1_weights[587][10] = -1;
        layer_1_weights[588][10] = 0;
        layer_1_weights[589][10] = -3;
        layer_1_weights[590][10] = -4;
        layer_1_weights[591][10] = -1;
        layer_1_weights[592][10] = 1;
        layer_1_weights[593][10] = -1;
        layer_1_weights[594][10] = 0;
        layer_1_weights[595][10] = -2;
        layer_1_weights[596][10] = 0;
        layer_1_weights[597][10] = -3;
        layer_1_weights[598][10] = -1;
        layer_1_weights[599][10] = -2;
        layer_1_weights[600][10] = -1;
        layer_1_weights[601][10] = 0;
        layer_1_weights[602][10] = -2;
        layer_1_weights[603][10] = 0;
        layer_1_weights[604][10] = 0;
        layer_1_weights[605][10] = -1;
        layer_1_weights[606][10] = -3;
        layer_1_weights[607][10] = -2;
        layer_1_weights[608][10] = -1;
        layer_1_weights[609][10] = 1;
        layer_1_weights[610][10] = -2;
        layer_1_weights[611][10] = -1;
        layer_1_weights[612][10] = 0;
        layer_1_weights[613][10] = -3;
        layer_1_weights[614][10] = 2;
        layer_1_weights[615][10] = 2;
        layer_1_weights[616][10] = 1;
        layer_1_weights[617][10] = 2;
        layer_1_weights[618][10] = -4;
        layer_1_weights[619][10] = -1;
        layer_1_weights[620][10] = 1;
        layer_1_weights[621][10] = 1;
        layer_1_weights[622][10] = 1;
        layer_1_weights[623][10] = 0;
        layer_1_weights[624][10] = -1;
        layer_1_weights[625][10] = -2;
        layer_1_weights[626][10] = -1;
        layer_1_weights[627][10] = 0;
        layer_1_weights[628][10] = 2;
        layer_1_weights[629][10] = 1;
        layer_1_weights[630][10] = 1;
        layer_1_weights[631][10] = 0;
        layer_1_weights[632][10] = 0;
        layer_1_weights[633][10] = -1;
        layer_1_weights[634][10] = -1;
        layer_1_weights[635][10] = -2;
        layer_1_weights[636][10] = 0;
        layer_1_weights[637][10] = 0;
        layer_1_weights[638][10] = 0;
        layer_1_weights[639][10] = 0;
        layer_1_weights[640][10] = -1;
        layer_1_weights[641][10] = -1;
        layer_1_weights[642][10] = 2;
        layer_1_weights[643][10] = 2;
        layer_1_weights[644][10] = 0;
        layer_1_weights[645][10] = 0;
        layer_1_weights[646][10] = -5;
        layer_1_weights[647][10] = -1;
        layer_1_weights[648][10] = -5;
        layer_1_weights[649][10] = 0;
        layer_1_weights[650][10] = 0;
        layer_1_weights[651][10] = 0;
        layer_1_weights[652][10] = 1;
        layer_1_weights[653][10] = 0;
        layer_1_weights[654][10] = 2;
        layer_1_weights[655][10] = 1;
        layer_1_weights[656][10] = 2;
        layer_1_weights[657][10] = 1;
        layer_1_weights[658][10] = 1;
        layer_1_weights[659][10] = 2;
        layer_1_weights[660][10] = 0;
        layer_1_weights[661][10] = 0;
        layer_1_weights[662][10] = -1;
        layer_1_weights[663][10] = -1;
        layer_1_weights[664][10] = 0;
        layer_1_weights[665][10] = 0;
        layer_1_weights[666][10] = 2;
        layer_1_weights[667][10] = 0;
        layer_1_weights[668][10] = 0;
        layer_1_weights[669][10] = 2;
        layer_1_weights[670][10] = 0;
        layer_1_weights[671][10] = 0;
        layer_1_weights[672][10] = 0;
        layer_1_weights[673][10] = 0;
        layer_1_weights[674][10] = 3;
        layer_1_weights[675][10] = 1;
        layer_1_weights[676][10] = 1;
        layer_1_weights[677][10] = 1;
        layer_1_weights[678][10] = -1;
        layer_1_weights[679][10] = 2;
        layer_1_weights[680][10] = 0;
        layer_1_weights[681][10] = 1;
        layer_1_weights[682][10] = 0;
        layer_1_weights[683][10] = 3;
        layer_1_weights[684][10] = 0;
        layer_1_weights[685][10] = 0;
        layer_1_weights[686][10] = 2;
        layer_1_weights[687][10] = -1;
        layer_1_weights[688][10] = 1;
        layer_1_weights[689][10] = -2;
        layer_1_weights[690][10] = 0;
        layer_1_weights[691][10] = -1;
        layer_1_weights[692][10] = 1;
        layer_1_weights[693][10] = 1;
        layer_1_weights[694][10] = -1;
        layer_1_weights[695][10] = -1;
        layer_1_weights[696][10] = -4;
        layer_1_weights[697][10] = -4;
        layer_1_weights[698][10] = -2;
        layer_1_weights[699][10] = 0;
        layer_1_weights[700][10] = 0;
        layer_1_weights[701][10] = 0;
        layer_1_weights[702][10] = 1;
        layer_1_weights[703][10] = 1;
        layer_1_weights[704][10] = 0;
        layer_1_weights[705][10] = 0;
        layer_1_weights[706][10] = 0;
        layer_1_weights[707][10] = -1;
        layer_1_weights[708][10] = 2;
        layer_1_weights[709][10] = 2;
        layer_1_weights[710][10] = 3;
        layer_1_weights[711][10] = 2;
        layer_1_weights[712][10] = -2;
        layer_1_weights[713][10] = -1;
        layer_1_weights[714][10] = -1;
        layer_1_weights[715][10] = 0;
        layer_1_weights[716][10] = -1;
        layer_1_weights[717][10] = -1;
        layer_1_weights[718][10] = -2;
        layer_1_weights[719][10] = 2;
        layer_1_weights[720][10] = 0;
        layer_1_weights[721][10] = 0;
        layer_1_weights[722][10] = 1;
        layer_1_weights[723][10] = 2;
        layer_1_weights[724][10] = -2;
        layer_1_weights[725][10] = -1;
        layer_1_weights[726][10] = -2;
        layer_1_weights[727][10] = -1;
        layer_1_weights[728][10] = 0;
        layer_1_weights[729][10] = 0;
        layer_1_weights[730][10] = 0;
        layer_1_weights[731][10] = 2;
        layer_1_weights[732][10] = -2;
        layer_1_weights[733][10] = -2;
        layer_1_weights[734][10] = -1;
        layer_1_weights[735][10] = 3;
        layer_1_weights[736][10] = 1;
        layer_1_weights[737][10] = 3;
        layer_1_weights[738][10] = -1;
        layer_1_weights[739][10] = 0;
        layer_1_weights[740][10] = 1;
        layer_1_weights[741][10] = 2;
        layer_1_weights[742][10] = 1;
        layer_1_weights[743][10] = 2;
        layer_1_weights[744][10] = 0;
        layer_1_weights[745][10] = 2;
        layer_1_weights[746][10] = 2;
        layer_1_weights[747][10] = 0;
        layer_1_weights[748][10] = 1;
        layer_1_weights[749][10] = 3;
        layer_1_weights[750][10] = 0;
        layer_1_weights[751][10] = 1;
        layer_1_weights[752][10] = 0;
        layer_1_weights[753][10] = 2;
        layer_1_weights[754][10] = 1;
        layer_1_weights[755][10] = 0;
        layer_1_weights[756][10] = 0;
        layer_1_weights[757][10] = 1;
        layer_1_weights[758][10] = 0;
        layer_1_weights[759][10] = 0;
        layer_1_weights[760][10] = 2;
        layer_1_weights[761][10] = 2;
        layer_1_weights[762][10] = 1;
        layer_1_weights[763][10] = 2;
        layer_1_weights[764][10] = 3;
        layer_1_weights[765][10] = 5;
        layer_1_weights[766][10] = 2;
        layer_1_weights[767][10] = 2;
        layer_1_weights[768][10] = 0;
        layer_1_weights[769][10] = 1;
        layer_1_weights[770][10] = 8;
        layer_1_weights[771][10] = 6;
        layer_1_weights[772][10] = 7;
        layer_1_weights[773][10] = 10;
        layer_1_weights[774][10] = 6;
        layer_1_weights[775][10] = 6;
        layer_1_weights[776][10] = 4;
        layer_1_weights[777][10] = 5;
        layer_1_weights[778][10] = 4;
        layer_1_weights[779][10] = 2;
        layer_1_weights[780][10] = 0;
        layer_1_weights[781][10] = 0;
        layer_1_weights[782][10] = 1;
        layer_1_weights[783][10] = 0;
        layer_1_weights[0][11] = 0;
        layer_1_weights[1][11] = -1;
        layer_1_weights[2][11] = 0;
        layer_1_weights[3][11] = 1;
        layer_1_weights[4][11] = 0;
        layer_1_weights[5][11] = 0;
        layer_1_weights[6][11] = 0;
        layer_1_weights[7][11] = 1;
        layer_1_weights[8][11] = 0;
        layer_1_weights[9][11] = 0;
        layer_1_weights[10][11] = 0;
        layer_1_weights[11][11] = 0;
        layer_1_weights[12][11] = 1;
        layer_1_weights[13][11] = 0;
        layer_1_weights[14][11] = -2;
        layer_1_weights[15][11] = 0;
        layer_1_weights[16][11] = 0;
        layer_1_weights[17][11] = 0;
        layer_1_weights[18][11] = 0;
        layer_1_weights[19][11] = 0;
        layer_1_weights[20][11] = 0;
        layer_1_weights[21][11] = 0;
        layer_1_weights[22][11] = 0;
        layer_1_weights[23][11] = 0;
        layer_1_weights[24][11] = -1;
        layer_1_weights[25][11] = 0;
        layer_1_weights[26][11] = -1;
        layer_1_weights[27][11] = 0;
        layer_1_weights[28][11] = 0;
        layer_1_weights[29][11] = 0;
        layer_1_weights[30][11] = 0;
        layer_1_weights[31][11] = 0;
        layer_1_weights[32][11] = 0;
        layer_1_weights[33][11] = 2;
        layer_1_weights[34][11] = 3;
        layer_1_weights[35][11] = 4;
        layer_1_weights[36][11] = 3;
        layer_1_weights[37][11] = 3;
        layer_1_weights[38][11] = 4;
        layer_1_weights[39][11] = -1;
        layer_1_weights[40][11] = 1;
        layer_1_weights[41][11] = 0;
        layer_1_weights[42][11] = -3;
        layer_1_weights[43][11] = -1;
        layer_1_weights[44][11] = 0;
        layer_1_weights[45][11] = 0;
        layer_1_weights[46][11] = 4;
        layer_1_weights[47][11] = 4;
        layer_1_weights[48][11] = 4;
        layer_1_weights[49][11] = 4;
        layer_1_weights[50][11] = 3;
        layer_1_weights[51][11] = 2;
        layer_1_weights[52][11] = 1;
        layer_1_weights[53][11] = 0;
        layer_1_weights[54][11] = 0;
        layer_1_weights[55][11] = 0;
        layer_1_weights[56][11] = -1;
        layer_1_weights[57][11] = -1;
        layer_1_weights[58][11] = 1;
        layer_1_weights[59][11] = 0;
        layer_1_weights[60][11] = 3;
        layer_1_weights[61][11] = 2;
        layer_1_weights[62][11] = 0;
        layer_1_weights[63][11] = 3;
        layer_1_weights[64][11] = 2;
        layer_1_weights[65][11] = 2;
        layer_1_weights[66][11] = 4;
        layer_1_weights[67][11] = 4;
        layer_1_weights[68][11] = 3;
        layer_1_weights[69][11] = -1;
        layer_1_weights[70][11] = -3;
        layer_1_weights[71][11] = -1;
        layer_1_weights[72][11] = -3;
        layer_1_weights[73][11] = 0;
        layer_1_weights[74][11] = -1;
        layer_1_weights[75][11] = -1;
        layer_1_weights[76][11] = 0;
        layer_1_weights[77][11] = 2;
        layer_1_weights[78][11] = 1;
        layer_1_weights[79][11] = 0;
        layer_1_weights[80][11] = 5;
        layer_1_weights[81][11] = 2;
        layer_1_weights[82][11] = -1;
        layer_1_weights[83][11] = 1;
        layer_1_weights[84][11] = 0;
        layer_1_weights[85][11] = 0;
        layer_1_weights[86][11] = -2;
        layer_1_weights[87][11] = 2;
        layer_1_weights[88][11] = -1;
        layer_1_weights[89][11] = 4;
        layer_1_weights[90][11] = 5;
        layer_1_weights[91][11] = 4;
        layer_1_weights[92][11] = 1;
        layer_1_weights[93][11] = 0;
        layer_1_weights[94][11] = 0;
        layer_1_weights[95][11] = 3;
        layer_1_weights[96][11] = -1;
        layer_1_weights[97][11] = -1;
        layer_1_weights[98][11] = 1;
        layer_1_weights[99][11] = -1;
        layer_1_weights[100][11] = 0;
        layer_1_weights[101][11] = 1;
        layer_1_weights[102][11] = -2;
        layer_1_weights[103][11] = -1;
        layer_1_weights[104][11] = -1;
        layer_1_weights[105][11] = -1;
        layer_1_weights[106][11] = -2;
        layer_1_weights[107][11] = 1;
        layer_1_weights[108][11] = -1;
        layer_1_weights[109][11] = 1;
        layer_1_weights[110][11] = 2;
        layer_1_weights[111][11] = -1;
        layer_1_weights[112][11] = 0;
        layer_1_weights[113][11] = 0;
        layer_1_weights[114][11] = -2;
        layer_1_weights[115][11] = -1;
        layer_1_weights[116][11] = 1;
        layer_1_weights[117][11] = 3;
        layer_1_weights[118][11] = 1;
        layer_1_weights[119][11] = -2;
        layer_1_weights[120][11] = -1;
        layer_1_weights[121][11] = -1;
        layer_1_weights[122][11] = 0;
        layer_1_weights[123][11] = -1;
        layer_1_weights[124][11] = -1;
        layer_1_weights[125][11] = -2;
        layer_1_weights[126][11] = -1;
        layer_1_weights[127][11] = -2;
        layer_1_weights[128][11] = 1;
        layer_1_weights[129][11] = -1;
        layer_1_weights[130][11] = 0;
        layer_1_weights[131][11] = 0;
        layer_1_weights[132][11] = 1;
        layer_1_weights[133][11] = 0;
        layer_1_weights[134][11] = 0;
        layer_1_weights[135][11] = -1;
        layer_1_weights[136][11] = -1;
        layer_1_weights[137][11] = 1;
        layer_1_weights[138][11] = -2;
        layer_1_weights[139][11] = -1;
        layer_1_weights[140][11] = -1;
        layer_1_weights[141][11] = 1;
        layer_1_weights[142][11] = 5;
        layer_1_weights[143][11] = -3;
        layer_1_weights[144][11] = 2;
        layer_1_weights[145][11] = 3;
        layer_1_weights[146][11] = 0;
        layer_1_weights[147][11] = 0;
        layer_1_weights[148][11] = -1;
        layer_1_weights[149][11] = -1;
        layer_1_weights[150][11] = -1;
        layer_1_weights[151][11] = -2;
        layer_1_weights[152][11] = -2;
        layer_1_weights[153][11] = 0;
        layer_1_weights[154][11] = 1;
        layer_1_weights[155][11] = -1;
        layer_1_weights[156][11] = 0;
        layer_1_weights[157][11] = -1;
        layer_1_weights[158][11] = 1;
        layer_1_weights[159][11] = -1;
        layer_1_weights[160][11] = 0;
        layer_1_weights[161][11] = -1;
        layer_1_weights[162][11] = -2;
        layer_1_weights[163][11] = 0;
        layer_1_weights[164][11] = 2;
        layer_1_weights[165][11] = -2;
        layer_1_weights[166][11] = 1;
        layer_1_weights[167][11] = -2;
        layer_1_weights[168][11] = 0;
        layer_1_weights[169][11] = 0;
        layer_1_weights[170][11] = -1;
        layer_1_weights[171][11] = -1;
        layer_1_weights[172][11] = 3;
        layer_1_weights[173][11] = 3;
        layer_1_weights[174][11] = 0;
        layer_1_weights[175][11] = 0;
        layer_1_weights[176][11] = 2;
        layer_1_weights[177][11] = 0;
        layer_1_weights[178][11] = -1;
        layer_1_weights[179][11] = 0;
        layer_1_weights[180][11] = -1;
        layer_1_weights[181][11] = 0;
        layer_1_weights[182][11] = -1;
        layer_1_weights[183][11] = 1;
        layer_1_weights[184][11] = -1;
        layer_1_weights[185][11] = 1;
        layer_1_weights[186][11] = -1;
        layer_1_weights[187][11] = 0;
        layer_1_weights[188][11] = -1;
        layer_1_weights[189][11] = -2;
        layer_1_weights[190][11] = 0;
        layer_1_weights[191][11] = -2;
        layer_1_weights[192][11] = -3;
        layer_1_weights[193][11] = -1;
        layer_1_weights[194][11] = 0;
        layer_1_weights[195][11] = 1;
        layer_1_weights[196][11] = -1;
        layer_1_weights[197][11] = -4;
        layer_1_weights[198][11] = 0;
        layer_1_weights[199][11] = -2;
        layer_1_weights[200][11] = 0;
        layer_1_weights[201][11] = 0;
        layer_1_weights[202][11] = -1;
        layer_1_weights[203][11] = 0;
        layer_1_weights[204][11] = -1;
        layer_1_weights[205][11] = 1;
        layer_1_weights[206][11] = -1;
        layer_1_weights[207][11] = 0;
        layer_1_weights[208][11] = -2;
        layer_1_weights[209][11] = 0;
        layer_1_weights[210][11] = -2;
        layer_1_weights[211][11] = 1;
        layer_1_weights[212][11] = 0;
        layer_1_weights[213][11] = 1;
        layer_1_weights[214][11] = 0;
        layer_1_weights[215][11] = 0;
        layer_1_weights[216][11] = -1;
        layer_1_weights[217][11] = 1;
        layer_1_weights[218][11] = -1;
        layer_1_weights[219][11] = -4;
        layer_1_weights[220][11] = 1;
        layer_1_weights[221][11] = 1;
        layer_1_weights[222][11] = 1;
        layer_1_weights[223][11] = 0;
        layer_1_weights[224][11] = -2;
        layer_1_weights[225][11] = 1;
        layer_1_weights[226][11] = 1;
        layer_1_weights[227][11] = -2;
        layer_1_weights[228][11] = -1;
        layer_1_weights[229][11] = -1;
        layer_1_weights[230][11] = 0;
        layer_1_weights[231][11] = -1;
        layer_1_weights[232][11] = -1;
        layer_1_weights[233][11] = -1;
        layer_1_weights[234][11] = -1;
        layer_1_weights[235][11] = -1;
        layer_1_weights[236][11] = -2;
        layer_1_weights[237][11] = 0;
        layer_1_weights[238][11] = -1;
        layer_1_weights[239][11] = 1;
        layer_1_weights[240][11] = 0;
        layer_1_weights[241][11] = 0;
        layer_1_weights[242][11] = 1;
        layer_1_weights[243][11] = 0;
        layer_1_weights[244][11] = 2;
        layer_1_weights[245][11] = 1;
        layer_1_weights[246][11] = -1;
        layer_1_weights[247][11] = 1;
        layer_1_weights[248][11] = -3;
        layer_1_weights[249][11] = -1;
        layer_1_weights[250][11] = 1;
        layer_1_weights[251][11] = -2;
        layer_1_weights[252][11] = -1;
        layer_1_weights[253][11] = -1;
        layer_1_weights[254][11] = -3;
        layer_1_weights[255][11] = 0;
        layer_1_weights[256][11] = -1;
        layer_1_weights[257][11] = -1;
        layer_1_weights[258][11] = 0;
        layer_1_weights[259][11] = 2;
        layer_1_weights[260][11] = 0;
        layer_1_weights[261][11] = 0;
        layer_1_weights[262][11] = 0;
        layer_1_weights[263][11] = 0;
        layer_1_weights[264][11] = 0;
        layer_1_weights[265][11] = -1;
        layer_1_weights[266][11] = -1;
        layer_1_weights[267][11] = -1;
        layer_1_weights[268][11] = -1;
        layer_1_weights[269][11] = -2;
        layer_1_weights[270][11] = 0;
        layer_1_weights[271][11] = -1;
        layer_1_weights[272][11] = 0;
        layer_1_weights[273][11] = -1;
        layer_1_weights[274][11] = -2;
        layer_1_weights[275][11] = -2;
        layer_1_weights[276][11] = -4;
        layer_1_weights[277][11] = -2;
        layer_1_weights[278][11] = -2;
        layer_1_weights[279][11] = -2;
        layer_1_weights[280][11] = -1;
        layer_1_weights[281][11] = -1;
        layer_1_weights[282][11] = -4;
        layer_1_weights[283][11] = 1;
        layer_1_weights[284][11] = -4;
        layer_1_weights[285][11] = 1;
        layer_1_weights[286][11] = 1;
        layer_1_weights[287][11] = 0;
        layer_1_weights[288][11] = 0;
        layer_1_weights[289][11] = 0;
        layer_1_weights[290][11] = -2;
        layer_1_weights[291][11] = -1;
        layer_1_weights[292][11] = -1;
        layer_1_weights[293][11] = -3;
        layer_1_weights[294][11] = -1;
        layer_1_weights[295][11] = -3;
        layer_1_weights[296][11] = 0;
        layer_1_weights[297][11] = -1;
        layer_1_weights[298][11] = 0;
        layer_1_weights[299][11] = 1;
        layer_1_weights[300][11] = 0;
        layer_1_weights[301][11] = 1;
        layer_1_weights[302][11] = -3;
        layer_1_weights[303][11] = -2;
        layer_1_weights[304][11] = -4;
        layer_1_weights[305][11] = 0;
        layer_1_weights[306][11] = -5;
        layer_1_weights[307][11] = -1;
        layer_1_weights[308][11] = -1;
        layer_1_weights[309][11] = -4;
        layer_1_weights[310][11] = 0;
        layer_1_weights[311][11] = -3;
        layer_1_weights[312][11] = -1;
        layer_1_weights[313][11] = 1;
        layer_1_weights[314][11] = 0;
        layer_1_weights[315][11] = 1;
        layer_1_weights[316][11] = 0;
        layer_1_weights[317][11] = 1;
        layer_1_weights[318][11] = 1;
        layer_1_weights[319][11] = -1;
        layer_1_weights[320][11] = -1;
        layer_1_weights[321][11] = -1;
        layer_1_weights[322][11] = -3;
        layer_1_weights[323][11] = -2;
        layer_1_weights[324][11] = -2;
        layer_1_weights[325][11] = -2;
        layer_1_weights[326][11] = -1;
        layer_1_weights[327][11] = 1;
        layer_1_weights[328][11] = 0;
        layer_1_weights[329][11] = 0;
        layer_1_weights[330][11] = 0;
        layer_1_weights[331][11] = 1;
        layer_1_weights[332][11] = -4;
        layer_1_weights[333][11] = -2;
        layer_1_weights[334][11] = -5;
        layer_1_weights[335][11] = -2;
        layer_1_weights[336][11] = -1;
        layer_1_weights[337][11] = -2;
        layer_1_weights[338][11] = -1;
        layer_1_weights[339][11] = -2;
        layer_1_weights[340][11] = 0;
        layer_1_weights[341][11] = -1;
        layer_1_weights[342][11] = 0;
        layer_1_weights[343][11] = -1;
        layer_1_weights[344][11] = 0;
        layer_1_weights[345][11] = -1;
        layer_1_weights[346][11] = -1;
        layer_1_weights[347][11] = 0;
        layer_1_weights[348][11] = 1;
        layer_1_weights[349][11] = -1;
        layer_1_weights[350][11] = 0;
        layer_1_weights[351][11] = -2;
        layer_1_weights[352][11] = 0;
        layer_1_weights[353][11] = -2;
        layer_1_weights[354][11] = 1;
        layer_1_weights[355][11] = 0;
        layer_1_weights[356][11] = 0;
        layer_1_weights[357][11] = 0;
        layer_1_weights[358][11] = 0;
        layer_1_weights[359][11] = 0;
        layer_1_weights[360][11] = -3;
        layer_1_weights[361][11] = -3;
        layer_1_weights[362][11] = -2;
        layer_1_weights[363][11] = -3;
        layer_1_weights[364][11] = 0;
        layer_1_weights[365][11] = 0;
        layer_1_weights[366][11] = -1;
        layer_1_weights[367][11] = -4;
        layer_1_weights[368][11] = -2;
        layer_1_weights[369][11] = -2;
        layer_1_weights[370][11] = 3;
        layer_1_weights[371][11] = 0;
        layer_1_weights[372][11] = 0;
        layer_1_weights[373][11] = -1;
        layer_1_weights[374][11] = 1;
        layer_1_weights[375][11] = -2;
        layer_1_weights[376][11] = 0;
        layer_1_weights[377][11] = 0;
        layer_1_weights[378][11] = 1;
        layer_1_weights[379][11] = 0;
        layer_1_weights[380][11] = -1;
        layer_1_weights[381][11] = -2;
        layer_1_weights[382][11] = -1;
        layer_1_weights[383][11] = 1;
        layer_1_weights[384][11] = 2;
        layer_1_weights[385][11] = 1;
        layer_1_weights[386][11] = 1;
        layer_1_weights[387][11] = 1;
        layer_1_weights[388][11] = 1;
        layer_1_weights[389][11] = -2;
        layer_1_weights[390][11] = 0;
        layer_1_weights[391][11] = -1;
        layer_1_weights[392][11] = -3;
        layer_1_weights[393][11] = 0;
        layer_1_weights[394][11] = -3;
        layer_1_weights[395][11] = 0;
        layer_1_weights[396][11] = 1;
        layer_1_weights[397][11] = 1;
        layer_1_weights[398][11] = 2;
        layer_1_weights[399][11] = 2;
        layer_1_weights[400][11] = 0;
        layer_1_weights[401][11] = 2;
        layer_1_weights[402][11] = 0;
        layer_1_weights[403][11] = 0;
        layer_1_weights[404][11] = 0;
        layer_1_weights[405][11] = -1;
        layer_1_weights[406][11] = 0;
        layer_1_weights[407][11] = -1;
        layer_1_weights[408][11] = 1;
        layer_1_weights[409][11] = -1;
        layer_1_weights[410][11] = 0;
        layer_1_weights[411][11] = 2;
        layer_1_weights[412][11] = 3;
        layer_1_weights[413][11] = 2;
        layer_1_weights[414][11] = 3;
        layer_1_weights[415][11] = 0;
        layer_1_weights[416][11] = 0;
        layer_1_weights[417][11] = -2;
        layer_1_weights[418][11] = -2;
        layer_1_weights[419][11] = 3;
        layer_1_weights[420][11] = -2;
        layer_1_weights[421][11] = -1;
        layer_1_weights[422][11] = -4;
        layer_1_weights[423][11] = -1;
        layer_1_weights[424][11] = 2;
        layer_1_weights[425][11] = 2;
        layer_1_weights[426][11] = 3;
        layer_1_weights[427][11] = 2;
        layer_1_weights[428][11] = 0;
        layer_1_weights[429][11] = 3;
        layer_1_weights[430][11] = 0;
        layer_1_weights[431][11] = 1;
        layer_1_weights[432][11] = 0;
        layer_1_weights[433][11] = 1;
        layer_1_weights[434][11] = 0;
        layer_1_weights[435][11] = 0;
        layer_1_weights[436][11] = 0;
        layer_1_weights[437][11] = 1;
        layer_1_weights[438][11] = 2;
        layer_1_weights[439][11] = 3;
        layer_1_weights[440][11] = 3;
        layer_1_weights[441][11] = 2;
        layer_1_weights[442][11] = 1;
        layer_1_weights[443][11] = 2;
        layer_1_weights[444][11] = -2;
        layer_1_weights[445][11] = 2;
        layer_1_weights[446][11] = -2;
        layer_1_weights[447][11] = 1;
        layer_1_weights[448][11] = 0;
        layer_1_weights[449][11] = -2;
        layer_1_weights[450][11] = 1;
        layer_1_weights[451][11] = -1;
        layer_1_weights[452][11] = 0;
        layer_1_weights[453][11] = 2;
        layer_1_weights[454][11] = 0;
        layer_1_weights[455][11] = 2;
        layer_1_weights[456][11] = 3;
        layer_1_weights[457][11] = 1;
        layer_1_weights[458][11] = 2;
        layer_1_weights[459][11] = 3;
        layer_1_weights[460][11] = 1;
        layer_1_weights[461][11] = 1;
        layer_1_weights[462][11] = 0;
        layer_1_weights[463][11] = 0;
        layer_1_weights[464][11] = 0;
        layer_1_weights[465][11] = 2;
        layer_1_weights[466][11] = 3;
        layer_1_weights[467][11] = 3;
        layer_1_weights[468][11] = 1;
        layer_1_weights[469][11] = 2;
        layer_1_weights[470][11] = 1;
        layer_1_weights[471][11] = 0;
        layer_1_weights[472][11] = -2;
        layer_1_weights[473][11] = 1;
        layer_1_weights[474][11] = 1;
        layer_1_weights[475][11] = 2;
        layer_1_weights[476][11] = 0;
        layer_1_weights[477][11] = -1;
        layer_1_weights[478][11] = 0;
        layer_1_weights[479][11] = -3;
        layer_1_weights[480][11] = -2;
        layer_1_weights[481][11] = -1;
        layer_1_weights[482][11] = 2;
        layer_1_weights[483][11] = 3;
        layer_1_weights[484][11] = 3;
        layer_1_weights[485][11] = 2;
        layer_1_weights[486][11] = 3;
        layer_1_weights[487][11] = 2;
        layer_1_weights[488][11] = 2;
        layer_1_weights[489][11] = 0;
        layer_1_weights[490][11] = 1;
        layer_1_weights[491][11] = 3;
        layer_1_weights[492][11] = 3;
        layer_1_weights[493][11] = 3;
        layer_1_weights[494][11] = 2;
        layer_1_weights[495][11] = 3;
        layer_1_weights[496][11] = 1;
        layer_1_weights[497][11] = 2;
        layer_1_weights[498][11] = 1;
        layer_1_weights[499][11] = -1;
        layer_1_weights[500][11] = -3;
        layer_1_weights[501][11] = 4;
        layer_1_weights[502][11] = -1;
        layer_1_weights[503][11] = -1;
        layer_1_weights[504][11] = 0;
        layer_1_weights[505][11] = 0;
        layer_1_weights[506][11] = -1;
        layer_1_weights[507][11] = 2;
        layer_1_weights[508][11] = 2;
        layer_1_weights[509][11] = 0;
        layer_1_weights[510][11] = 1;
        layer_1_weights[511][11] = 3;
        layer_1_weights[512][11] = 1;
        layer_1_weights[513][11] = 1;
        layer_1_weights[514][11] = 1;
        layer_1_weights[515][11] = 2;
        layer_1_weights[516][11] = 1;
        layer_1_weights[517][11] = 2;
        layer_1_weights[518][11] = 2;
        layer_1_weights[519][11] = 3;
        layer_1_weights[520][11] = 4;
        layer_1_weights[521][11] = 4;
        layer_1_weights[522][11] = 4;
        layer_1_weights[523][11] = 2;
        layer_1_weights[524][11] = 0;
        layer_1_weights[525][11] = 0;
        layer_1_weights[526][11] = 2;
        layer_1_weights[527][11] = -1;
        layer_1_weights[528][11] = -2;
        layer_1_weights[529][11] = 0;
        layer_1_weights[530][11] = 0;
        layer_1_weights[531][11] = 1;
        layer_1_weights[532][11] = 0;
        layer_1_weights[533][11] = -3;
        layer_1_weights[534][11] = -1;
        layer_1_weights[535][11] = 1;
        layer_1_weights[536][11] = 0;
        layer_1_weights[537][11] = -1;
        layer_1_weights[538][11] = -1;
        layer_1_weights[539][11] = -1;
        layer_1_weights[540][11] = 0;
        layer_1_weights[541][11] = 0;
        layer_1_weights[542][11] = 0;
        layer_1_weights[543][11] = 3;
        layer_1_weights[544][11] = 0;
        layer_1_weights[545][11] = 2;
        layer_1_weights[546][11] = 2;
        layer_1_weights[547][11] = 3;
        layer_1_weights[548][11] = 3;
        layer_1_weights[549][11] = 2;
        layer_1_weights[550][11] = 2;
        layer_1_weights[551][11] = 2;
        layer_1_weights[552][11] = 2;
        layer_1_weights[553][11] = 0;
        layer_1_weights[554][11] = -1;
        layer_1_weights[555][11] = -1;
        layer_1_weights[556][11] = 2;
        layer_1_weights[557][11] = -2;
        layer_1_weights[558][11] = 3;
        layer_1_weights[559][11] = -1;
        layer_1_weights[560][11] = 1;
        layer_1_weights[561][11] = -2;
        layer_1_weights[562][11] = 4;
        layer_1_weights[563][11] = 2;
        layer_1_weights[564][11] = -1;
        layer_1_weights[565][11] = -1;
        layer_1_weights[566][11] = -2;
        layer_1_weights[567][11] = -3;
        layer_1_weights[568][11] = 0;
        layer_1_weights[569][11] = -1;
        layer_1_weights[570][11] = 0;
        layer_1_weights[571][11] = 0;
        layer_1_weights[572][11] = 0;
        layer_1_weights[573][11] = 0;
        layer_1_weights[574][11] = 1;
        layer_1_weights[575][11] = 1;
        layer_1_weights[576][11] = 1;
        layer_1_weights[577][11] = 0;
        layer_1_weights[578][11] = 1;
        layer_1_weights[579][11] = 0;
        layer_1_weights[580][11] = 0;
        layer_1_weights[581][11] = -1;
        layer_1_weights[582][11] = 1;
        layer_1_weights[583][11] = -1;
        layer_1_weights[584][11] = 0;
        layer_1_weights[585][11] = 0;
        layer_1_weights[586][11] = 4;
        layer_1_weights[587][11] = 0;
        layer_1_weights[588][11] = 0;
        layer_1_weights[589][11] = 0;
        layer_1_weights[590][11] = 2;
        layer_1_weights[591][11] = 1;
        layer_1_weights[592][11] = 0;
        layer_1_weights[593][11] = 0;
        layer_1_weights[594][11] = -3;
        layer_1_weights[595][11] = 1;
        layer_1_weights[596][11] = -1;
        layer_1_weights[597][11] = -2;
        layer_1_weights[598][11] = -1;
        layer_1_weights[599][11] = -2;
        layer_1_weights[600][11] = 1;
        layer_1_weights[601][11] = 0;
        layer_1_weights[602][11] = 1;
        layer_1_weights[603][11] = 0;
        layer_1_weights[604][11] = 1;
        layer_1_weights[605][11] = 0;
        layer_1_weights[606][11] = 1;
        layer_1_weights[607][11] = 1;
        layer_1_weights[608][11] = -2;
        layer_1_weights[609][11] = -2;
        layer_1_weights[610][11] = -1;
        layer_1_weights[611][11] = -1;
        layer_1_weights[612][11] = 1;
        layer_1_weights[613][11] = -1;
        layer_1_weights[614][11] = 1;
        layer_1_weights[615][11] = 0;
        layer_1_weights[616][11] = 1;
        layer_1_weights[617][11] = 0;
        layer_1_weights[618][11] = 1;
        layer_1_weights[619][11] = -1;
        layer_1_weights[620][11] = 0;
        layer_1_weights[621][11] = -1;
        layer_1_weights[622][11] = -1;
        layer_1_weights[623][11] = -1;
        layer_1_weights[624][11] = -2;
        layer_1_weights[625][11] = 0;
        layer_1_weights[626][11] = 0;
        layer_1_weights[627][11] = -1;
        layer_1_weights[628][11] = 1;
        layer_1_weights[629][11] = 0;
        layer_1_weights[630][11] = -3;
        layer_1_weights[631][11] = -2;
        layer_1_weights[632][11] = 0;
        layer_1_weights[633][11] = -2;
        layer_1_weights[634][11] = -3;
        layer_1_weights[635][11] = -1;
        layer_1_weights[636][11] = -3;
        layer_1_weights[637][11] = -1;
        layer_1_weights[638][11] = -1;
        layer_1_weights[639][11] = -1;
        layer_1_weights[640][11] = -1;
        layer_1_weights[641][11] = -2;
        layer_1_weights[642][11] = -1;
        layer_1_weights[643][11] = 0;
        layer_1_weights[644][11] = 1;
        layer_1_weights[645][11] = 0;
        layer_1_weights[646][11] = 0;
        layer_1_weights[647][11] = 0;
        layer_1_weights[648][11] = 2;
        layer_1_weights[649][11] = 1;
        layer_1_weights[650][11] = -1;
        layer_1_weights[651][11] = -1;
        layer_1_weights[652][11] = -2;
        layer_1_weights[653][11] = -1;
        layer_1_weights[654][11] = -1;
        layer_1_weights[655][11] = -1;
        layer_1_weights[656][11] = -1;
        layer_1_weights[657][11] = -1;
        layer_1_weights[658][11] = -2;
        layer_1_weights[659][11] = -1;
        layer_1_weights[660][11] = -1;
        layer_1_weights[661][11] = -2;
        layer_1_weights[662][11] = -3;
        layer_1_weights[663][11] = -1;
        layer_1_weights[664][11] = 0;
        layer_1_weights[665][11] = -2;
        layer_1_weights[666][11] = -1;
        layer_1_weights[667][11] = -1;
        layer_1_weights[668][11] = 0;
        layer_1_weights[669][11] = -3;
        layer_1_weights[670][11] = -3;
        layer_1_weights[671][11] = 0;
        layer_1_weights[672][11] = 0;
        layer_1_weights[673][11] = 0;
        layer_1_weights[674][11] = 1;
        layer_1_weights[675][11] = -1;
        layer_1_weights[676][11] = -1;
        layer_1_weights[677][11] = 4;
        layer_1_weights[678][11] = 0;
        layer_1_weights[679][11] = 2;
        layer_1_weights[680][11] = 2;
        layer_1_weights[681][11] = 0;
        layer_1_weights[682][11] = 0;
        layer_1_weights[683][11] = 1;
        layer_1_weights[684][11] = -1;
        layer_1_weights[685][11] = -2;
        layer_1_weights[686][11] = -2;
        layer_1_weights[687][11] = -1;
        layer_1_weights[688][11] = -2;
        layer_1_weights[689][11] = -1;
        layer_1_weights[690][11] = -2;
        layer_1_weights[691][11] = -4;
        layer_1_weights[692][11] = -1;
        layer_1_weights[693][11] = -1;
        layer_1_weights[694][11] = -2;
        layer_1_weights[695][11] = 1;
        layer_1_weights[696][11] = -1;
        layer_1_weights[697][11] = 2;
        layer_1_weights[698][11] = 0;
        layer_1_weights[699][11] = 0;
        layer_1_weights[700][11] = 0;
        layer_1_weights[701][11] = 0;
        layer_1_weights[702][11] = 2;
        layer_1_weights[703][11] = -1;
        layer_1_weights[704][11] = 0;
        layer_1_weights[705][11] = 3;
        layer_1_weights[706][11] = 1;
        layer_1_weights[707][11] = 0;
        layer_1_weights[708][11] = 1;
        layer_1_weights[709][11] = 0;
        layer_1_weights[710][11] = -2;
        layer_1_weights[711][11] = 0;
        layer_1_weights[712][11] = 0;
        layer_1_weights[713][11] = 1;
        layer_1_weights[714][11] = -1;
        layer_1_weights[715][11] = 0;
        layer_1_weights[716][11] = -2;
        layer_1_weights[717][11] = -2;
        layer_1_weights[718][11] = -2;
        layer_1_weights[719][11] = 3;
        layer_1_weights[720][11] = 0;
        layer_1_weights[721][11] = 3;
        layer_1_weights[722][11] = 1;
        layer_1_weights[723][11] = 0;
        layer_1_weights[724][11] = -3;
        layer_1_weights[725][11] = 2;
        layer_1_weights[726][11] = 0;
        layer_1_weights[727][11] = 0;
        layer_1_weights[728][11] = 0;
        layer_1_weights[729][11] = 0;
        layer_1_weights[730][11] = 0;
        layer_1_weights[731][11] = 1;
        layer_1_weights[732][11] = 2;
        layer_1_weights[733][11] = 4;
        layer_1_weights[734][11] = 6;
        layer_1_weights[735][11] = 5;
        layer_1_weights[736][11] = 4;
        layer_1_weights[737][11] = 4;
        layer_1_weights[738][11] = 2;
        layer_1_weights[739][11] = 0;
        layer_1_weights[740][11] = 1;
        layer_1_weights[741][11] = 2;
        layer_1_weights[742][11] = 3;
        layer_1_weights[743][11] = 3;
        layer_1_weights[744][11] = -1;
        layer_1_weights[745][11] = 0;
        layer_1_weights[746][11] = -1;
        layer_1_weights[747][11] = -1;
        layer_1_weights[748][11] = 2;
        layer_1_weights[749][11] = 3;
        layer_1_weights[750][11] = -1;
        layer_1_weights[751][11] = 3;
        layer_1_weights[752][11] = -1;
        layer_1_weights[753][11] = -1;
        layer_1_weights[754][11] = 0;
        layer_1_weights[755][11] = 0;
        layer_1_weights[756][11] = -1;
        layer_1_weights[757][11] = -1;
        layer_1_weights[758][11] = 0;
        layer_1_weights[759][11] = 0;
        layer_1_weights[760][11] = -2;
        layer_1_weights[761][11] = -4;
        layer_1_weights[762][11] = 2;
        layer_1_weights[763][11] = 1;
        layer_1_weights[764][11] = 2;
        layer_1_weights[765][11] = 2;
        layer_1_weights[766][11] = 1;
        layer_1_weights[767][11] = 0;
        layer_1_weights[768][11] = 0;
        layer_1_weights[769][11] = -1;
        layer_1_weights[770][11] = -1;
        layer_1_weights[771][11] = 0;
        layer_1_weights[772][11] = 0;
        layer_1_weights[773][11] = -2;
        layer_1_weights[774][11] = 1;
        layer_1_weights[775][11] = 1;
        layer_1_weights[776][11] = 2;
        layer_1_weights[777][11] = -1;
        layer_1_weights[778][11] = 0;
        layer_1_weights[779][11] = -3;
        layer_1_weights[780][11] = 0;
        layer_1_weights[781][11] = 0;
        layer_1_weights[782][11] = 0;
        layer_1_weights[783][11] = -1;
        layer_1_weights[0][12] = 0;
        layer_1_weights[1][12] = 0;
        layer_1_weights[2][12] = 0;
        layer_1_weights[3][12] = 0;
        layer_1_weights[4][12] = 0;
        layer_1_weights[5][12] = 0;
        layer_1_weights[6][12] = 0;
        layer_1_weights[7][12] = -1;
        layer_1_weights[8][12] = -1;
        layer_1_weights[9][12] = 0;
        layer_1_weights[10][12] = 0;
        layer_1_weights[11][12] = 0;
        layer_1_weights[12][12] = 1;
        layer_1_weights[13][12] = 2;
        layer_1_weights[14][12] = -1;
        layer_1_weights[15][12] = -1;
        layer_1_weights[16][12] = 1;
        layer_1_weights[17][12] = 0;
        layer_1_weights[18][12] = 0;
        layer_1_weights[19][12] = 0;
        layer_1_weights[20][12] = 1;
        layer_1_weights[21][12] = 0;
        layer_1_weights[22][12] = 0;
        layer_1_weights[23][12] = 0;
        layer_1_weights[24][12] = 1;
        layer_1_weights[25][12] = 0;
        layer_1_weights[26][12] = 0;
        layer_1_weights[27][12] = 0;
        layer_1_weights[28][12] = 0;
        layer_1_weights[29][12] = 0;
        layer_1_weights[30][12] = 0;
        layer_1_weights[31][12] = 0;
        layer_1_weights[32][12] = 0;
        layer_1_weights[33][12] = 2;
        layer_1_weights[34][12] = 1;
        layer_1_weights[35][12] = 2;
        layer_1_weights[36][12] = 0;
        layer_1_weights[37][12] = 2;
        layer_1_weights[38][12] = 4;
        layer_1_weights[39][12] = 0;
        layer_1_weights[40][12] = 1;
        layer_1_weights[41][12] = 2;
        layer_1_weights[42][12] = 3;
        layer_1_weights[43][12] = -1;
        layer_1_weights[44][12] = 0;
        layer_1_weights[45][12] = 1;
        layer_1_weights[46][12] = 5;
        layer_1_weights[47][12] = 5;
        layer_1_weights[48][12] = 5;
        layer_1_weights[49][12] = 5;
        layer_1_weights[50][12] = 4;
        layer_1_weights[51][12] = 2;
        layer_1_weights[52][12] = 0;
        layer_1_weights[53][12] = 0;
        layer_1_weights[54][12] = 0;
        layer_1_weights[55][12] = 0;
        layer_1_weights[56][12] = 1;
        layer_1_weights[57][12] = 0;
        layer_1_weights[58][12] = 1;
        layer_1_weights[59][12] = 0;
        layer_1_weights[60][12] = 3;
        layer_1_weights[61][12] = 1;
        layer_1_weights[62][12] = 2;
        layer_1_weights[63][12] = 0;
        layer_1_weights[64][12] = -2;
        layer_1_weights[65][12] = -2;
        layer_1_weights[66][12] = -1;
        layer_1_weights[67][12] = 1;
        layer_1_weights[68][12] = 1;
        layer_1_weights[69][12] = 2;
        layer_1_weights[70][12] = 1;
        layer_1_weights[71][12] = 3;
        layer_1_weights[72][12] = 2;
        layer_1_weights[73][12] = 3;
        layer_1_weights[74][12] = 3;
        layer_1_weights[75][12] = 2;
        layer_1_weights[76][12] = 4;
        layer_1_weights[77][12] = 2;
        layer_1_weights[78][12] = 7;
        layer_1_weights[79][12] = 3;
        layer_1_weights[80][12] = 0;
        layer_1_weights[81][12] = 0;
        layer_1_weights[82][12] = 0;
        layer_1_weights[83][12] = 0;
        layer_1_weights[84][12] = 0;
        layer_1_weights[85][12] = 0;
        layer_1_weights[86][12] = -2;
        layer_1_weights[87][12] = 3;
        layer_1_weights[88][12] = 3;
        layer_1_weights[89][12] = -3;
        layer_1_weights[90][12] = -1;
        layer_1_weights[91][12] = -1;
        layer_1_weights[92][12] = -5;
        layer_1_weights[93][12] = -7;
        layer_1_weights[94][12] = -4;
        layer_1_weights[95][12] = -2;
        layer_1_weights[96][12] = -1;
        layer_1_weights[97][12] = -1;
        layer_1_weights[98][12] = -2;
        layer_1_weights[99][12] = -1;
        layer_1_weights[100][12] = 2;
        layer_1_weights[101][12] = 0;
        layer_1_weights[102][12] = 5;
        layer_1_weights[103][12] = 4;
        layer_1_weights[104][12] = 1;
        layer_1_weights[105][12] = 2;
        layer_1_weights[106][12] = 3;
        layer_1_weights[107][12] = 6;
        layer_1_weights[108][12] = 3;
        layer_1_weights[109][12] = 1;
        layer_1_weights[110][12] = 2;
        layer_1_weights[111][12] = 0;
        layer_1_weights[112][12] = 0;
        layer_1_weights[113][12] = 0;
        layer_1_weights[114][12] = -4;
        layer_1_weights[115][12] = 1;
        layer_1_weights[116][12] = -2;
        layer_1_weights[117][12] = -4;
        layer_1_weights[118][12] = -5;
        layer_1_weights[119][12] = -4;
        layer_1_weights[120][12] = -4;
        layer_1_weights[121][12] = -1;
        layer_1_weights[122][12] = -1;
        layer_1_weights[123][12] = 0;
        layer_1_weights[124][12] = -2;
        layer_1_weights[125][12] = -1;
        layer_1_weights[126][12] = -1;
        layer_1_weights[127][12] = 0;
        layer_1_weights[128][12] = 0;
        layer_1_weights[129][12] = 0;
        layer_1_weights[130][12] = 0;
        layer_1_weights[131][12] = 0;
        layer_1_weights[132][12] = 1;
        layer_1_weights[133][12] = 0;
        layer_1_weights[134][12] = 1;
        layer_1_weights[135][12] = 3;
        layer_1_weights[136][12] = 2;
        layer_1_weights[137][12] = 2;
        layer_1_weights[138][12] = 4;
        layer_1_weights[139][12] = 3;
        layer_1_weights[140][12] = -1;
        layer_1_weights[141][12] = 1;
        layer_1_weights[142][12] = 4;
        layer_1_weights[143][12] = 1;
        layer_1_weights[144][12] = -2;
        layer_1_weights[145][12] = -4;
        layer_1_weights[146][12] = -3;
        layer_1_weights[147][12] = -2;
        layer_1_weights[148][12] = -3;
        layer_1_weights[149][12] = -1;
        layer_1_weights[150][12] = -1;
        layer_1_weights[151][12] = 0;
        layer_1_weights[152][12] = 0;
        layer_1_weights[153][12] = -1;
        layer_1_weights[154][12] = -1;
        layer_1_weights[155][12] = -1;
        layer_1_weights[156][12] = -2;
        layer_1_weights[157][12] = -1;
        layer_1_weights[158][12] = 0;
        layer_1_weights[159][12] = 0;
        layer_1_weights[160][12] = 2;
        layer_1_weights[161][12] = 0;
        layer_1_weights[162][12] = 0;
        layer_1_weights[163][12] = 1;
        layer_1_weights[164][12] = 1;
        layer_1_weights[165][12] = 2;
        layer_1_weights[166][12] = 7;
        layer_1_weights[167][12] = 3;
        layer_1_weights[168][12] = 0;
        layer_1_weights[169][12] = 0;
        layer_1_weights[170][12] = -1;
        layer_1_weights[171][12] = -6;
        layer_1_weights[172][12] = -2;
        layer_1_weights[173][12] = -2;
        layer_1_weights[174][12] = -3;
        layer_1_weights[175][12] = -2;
        layer_1_weights[176][12] = -2;
        layer_1_weights[177][12] = -2;
        layer_1_weights[178][12] = -1;
        layer_1_weights[179][12] = 0;
        layer_1_weights[180][12] = 0;
        layer_1_weights[181][12] = 1;
        layer_1_weights[182][12] = 1;
        layer_1_weights[183][12] = 2;
        layer_1_weights[184][12] = 1;
        layer_1_weights[185][12] = 1;
        layer_1_weights[186][12] = 0;
        layer_1_weights[187][12] = 0;
        layer_1_weights[188][12] = 1;
        layer_1_weights[189][12] = 0;
        layer_1_weights[190][12] = 1;
        layer_1_weights[191][12] = 1;
        layer_1_weights[192][12] = 3;
        layer_1_weights[193][12] = 8;
        layer_1_weights[194][12] = 5;
        layer_1_weights[195][12] = 2;
        layer_1_weights[196][12] = 1;
        layer_1_weights[197][12] = -4;
        layer_1_weights[198][12] = 1;
        layer_1_weights[199][12] = -3;
        layer_1_weights[200][12] = -3;
        layer_1_weights[201][12] = -3;
        layer_1_weights[202][12] = -3;
        layer_1_weights[203][12] = 0;
        layer_1_weights[204][12] = 0;
        layer_1_weights[205][12] = -1;
        layer_1_weights[206][12] = 0;
        layer_1_weights[207][12] = -1;
        layer_1_weights[208][12] = -1;
        layer_1_weights[209][12] = 1;
        layer_1_weights[210][12] = 1;
        layer_1_weights[211][12] = 2;
        layer_1_weights[212][12] = 2;
        layer_1_weights[213][12] = 1;
        layer_1_weights[214][12] = 1;
        layer_1_weights[215][12] = 1;
        layer_1_weights[216][12] = 1;
        layer_1_weights[217][12] = 1;
        layer_1_weights[218][12] = 3;
        layer_1_weights[219][12] = 2;
        layer_1_weights[220][12] = 3;
        layer_1_weights[221][12] = 4;
        layer_1_weights[222][12] = 2;
        layer_1_weights[223][12] = 4;
        layer_1_weights[224][12] = 2;
        layer_1_weights[225][12] = -4;
        layer_1_weights[226][12] = -3;
        layer_1_weights[227][12] = -2;
        layer_1_weights[228][12] = -3;
        layer_1_weights[229][12] = -1;
        layer_1_weights[230][12] = -1;
        layer_1_weights[231][12] = 1;
        layer_1_weights[232][12] = 0;
        layer_1_weights[233][12] = 0;
        layer_1_weights[234][12] = 0;
        layer_1_weights[235][12] = 1;
        layer_1_weights[236][12] = 0;
        layer_1_weights[237][12] = 1;
        layer_1_weights[238][12] = 0;
        layer_1_weights[239][12] = 1;
        layer_1_weights[240][12] = 1;
        layer_1_weights[241][12] = 0;
        layer_1_weights[242][12] = 0;
        layer_1_weights[243][12] = -1;
        layer_1_weights[244][12] = -1;
        layer_1_weights[245][12] = 0;
        layer_1_weights[246][12] = 0;
        layer_1_weights[247][12] = 1;
        layer_1_weights[248][12] = 5;
        layer_1_weights[249][12] = 7;
        layer_1_weights[250][12] = 5;
        layer_1_weights[251][12] = 3;
        layer_1_weights[252][12] = 0;
        layer_1_weights[253][12] = -2;
        layer_1_weights[254][12] = -3;
        layer_1_weights[255][12] = -4;
        layer_1_weights[256][12] = -4;
        layer_1_weights[257][12] = -3;
        layer_1_weights[258][12] = 0;
        layer_1_weights[259][12] = 0;
        layer_1_weights[260][12] = 0;
        layer_1_weights[261][12] = 0;
        layer_1_weights[262][12] = 0;
        layer_1_weights[263][12] = 0;
        layer_1_weights[264][12] = 0;
        layer_1_weights[265][12] = 0;
        layer_1_weights[266][12] = 0;
        layer_1_weights[267][12] = -2;
        layer_1_weights[268][12] = -2;
        layer_1_weights[269][12] = -2;
        layer_1_weights[270][12] = -2;
        layer_1_weights[271][12] = -2;
        layer_1_weights[272][12] = -2;
        layer_1_weights[273][12] = 0;
        layer_1_weights[274][12] = -2;
        layer_1_weights[275][12] = -1;
        layer_1_weights[276][12] = 5;
        layer_1_weights[277][12] = 3;
        layer_1_weights[278][12] = 2;
        layer_1_weights[279][12] = -3;
        layer_1_weights[280][12] = -1;
        layer_1_weights[281][12] = 1;
        layer_1_weights[282][12] = -4;
        layer_1_weights[283][12] = -6;
        layer_1_weights[284][12] = -4;
        layer_1_weights[285][12] = -4;
        layer_1_weights[286][12] = -3;
        layer_1_weights[287][12] = 1;
        layer_1_weights[288][12] = 1;
        layer_1_weights[289][12] = 2;
        layer_1_weights[290][12] = 2;
        layer_1_weights[291][12] = 1;
        layer_1_weights[292][12] = -1;
        layer_1_weights[293][12] = 0;
        layer_1_weights[294][12] = -1;
        layer_1_weights[295][12] = -1;
        layer_1_weights[296][12] = -3;
        layer_1_weights[297][12] = -2;
        layer_1_weights[298][12] = -3;
        layer_1_weights[299][12] = -2;
        layer_1_weights[300][12] = -2;
        layer_1_weights[301][12] = -1;
        layer_1_weights[302][12] = -2;
        layer_1_weights[303][12] = 0;
        layer_1_weights[304][12] = 5;
        layer_1_weights[305][12] = 3;
        layer_1_weights[306][12] = 2;
        layer_1_weights[307][12] = -3;
        layer_1_weights[308][12] = 0;
        layer_1_weights[309][12] = 0;
        layer_1_weights[310][12] = 0;
        layer_1_weights[311][12] = -5;
        layer_1_weights[312][12] = -3;
        layer_1_weights[313][12] = 1;
        layer_1_weights[314][12] = -1;
        layer_1_weights[315][12] = 0;
        layer_1_weights[316][12] = 1;
        layer_1_weights[317][12] = 1;
        layer_1_weights[318][12] = 2;
        layer_1_weights[319][12] = 0;
        layer_1_weights[320][12] = 2;
        layer_1_weights[321][12] = 2;
        layer_1_weights[322][12] = 2;
        layer_1_weights[323][12] = 0;
        layer_1_weights[324][12] = -2;
        layer_1_weights[325][12] = -1;
        layer_1_weights[326][12] = -1;
        layer_1_weights[327][12] = -1;
        layer_1_weights[328][12] = -1;
        layer_1_weights[329][12] = -2;
        layer_1_weights[330][12] = -2;
        layer_1_weights[331][12] = 1;
        layer_1_weights[332][12] = 2;
        layer_1_weights[333][12] = 1;
        layer_1_weights[334][12] = 5;
        layer_1_weights[335][12] = 0;
        layer_1_weights[336][12] = -1;
        layer_1_weights[337][12] = -1;
        layer_1_weights[338][12] = -2;
        layer_1_weights[339][12] = -4;
        layer_1_weights[340][12] = -4;
        layer_1_weights[341][12] = -2;
        layer_1_weights[342][12] = 1;
        layer_1_weights[343][12] = 0;
        layer_1_weights[344][12] = 2;
        layer_1_weights[345][12] = 2;
        layer_1_weights[346][12] = 1;
        layer_1_weights[347][12] = 1;
        layer_1_weights[348][12] = 3;
        layer_1_weights[349][12] = 3;
        layer_1_weights[350][12] = 2;
        layer_1_weights[351][12] = 2;
        layer_1_weights[352][12] = 1;
        layer_1_weights[353][12] = 1;
        layer_1_weights[354][12] = 1;
        layer_1_weights[355][12] = -1;
        layer_1_weights[356][12] = 0;
        layer_1_weights[357][12] = 1;
        layer_1_weights[358][12] = -1;
        layer_1_weights[359][12] = 2;
        layer_1_weights[360][12] = 0;
        layer_1_weights[361][12] = -4;
        layer_1_weights[362][12] = -2;
        layer_1_weights[363][12] = -3;
        layer_1_weights[364][12] = 1;
        layer_1_weights[365][12] = -1;
        layer_1_weights[366][12] = -1;
        layer_1_weights[367][12] = -5;
        layer_1_weights[368][12] = -4;
        layer_1_weights[369][12] = -3;
        layer_1_weights[370][12] = 0;
        layer_1_weights[371][12] = -1;
        layer_1_weights[372][12] = 2;
        layer_1_weights[373][12] = 1;
        layer_1_weights[374][12] = 1;
        layer_1_weights[375][12] = 2;
        layer_1_weights[376][12] = 1;
        layer_1_weights[377][12] = 2;
        layer_1_weights[378][12] = 3;
        layer_1_weights[379][12] = 2;
        layer_1_weights[380][12] = 0;
        layer_1_weights[381][12] = 0;
        layer_1_weights[382][12] = 0;
        layer_1_weights[383][12] = 1;
        layer_1_weights[384][12] = 1;
        layer_1_weights[385][12] = 0;
        layer_1_weights[386][12] = 1;
        layer_1_weights[387][12] = -4;
        layer_1_weights[388][12] = -6;
        layer_1_weights[389][12] = -8;
        layer_1_weights[390][12] = -5;
        layer_1_weights[391][12] = 1;
        layer_1_weights[392][12] = 2;
        layer_1_weights[393][12] = 0;
        layer_1_weights[394][12] = -1;
        layer_1_weights[395][12] = -4;
        layer_1_weights[396][12] = -2;
        layer_1_weights[397][12] = -3;
        layer_1_weights[398][12] = 0;
        layer_1_weights[399][12] = 0;
        layer_1_weights[400][12] = 1;
        layer_1_weights[401][12] = 1;
        layer_1_weights[402][12] = 0;
        layer_1_weights[403][12] = 2;
        layer_1_weights[404][12] = 2;
        layer_1_weights[405][12] = 2;
        layer_1_weights[406][12] = 1;
        layer_1_weights[407][12] = 1;
        layer_1_weights[408][12] = 0;
        layer_1_weights[409][12] = 1;
        layer_1_weights[410][12] = -2;
        layer_1_weights[411][12] = -1;
        layer_1_weights[412][12] = 0;
        layer_1_weights[413][12] = 1;
        layer_1_weights[414][12] = 0;
        layer_1_weights[415][12] = 0;
        layer_1_weights[416][12] = -7;
        layer_1_weights[417][12] = -6;
        layer_1_weights[418][12] = -5;
        layer_1_weights[419][12] = -1;
        layer_1_weights[420][12] = 2;
        layer_1_weights[421][12] = 0;
        layer_1_weights[422][12] = -3;
        layer_1_weights[423][12] = -3;
        layer_1_weights[424][12] = -1;
        layer_1_weights[425][12] = -1;
        layer_1_weights[426][12] = 1;
        layer_1_weights[427][12] = -1;
        layer_1_weights[428][12] = 0;
        layer_1_weights[429][12] = 0;
        layer_1_weights[430][12] = 1;
        layer_1_weights[431][12] = 0;
        layer_1_weights[432][12] = 2;
        layer_1_weights[433][12] = 2;
        layer_1_weights[434][12] = 1;
        layer_1_weights[435][12] = -1;
        layer_1_weights[436][12] = 0;
        layer_1_weights[437][12] = -1;
        layer_1_weights[438][12] = -1;
        layer_1_weights[439][12] = -1;
        layer_1_weights[440][12] = -1;
        layer_1_weights[441][12] = 0;
        layer_1_weights[442][12] = -1;
        layer_1_weights[443][12] = -2;
        layer_1_weights[444][12] = -3;
        layer_1_weights[445][12] = -5;
        layer_1_weights[446][12] = -5;
        layer_1_weights[447][12] = -2;
        layer_1_weights[448][12] = -3;
        layer_1_weights[449][12] = -1;
        layer_1_weights[450][12] = -4;
        layer_1_weights[451][12] = -4;
        layer_1_weights[452][12] = -3;
        layer_1_weights[453][12] = -4;
        layer_1_weights[454][12] = -2;
        layer_1_weights[455][12] = -1;
        layer_1_weights[456][12] = -1;
        layer_1_weights[457][12] = -1;
        layer_1_weights[458][12] = 0;
        layer_1_weights[459][12] = 2;
        layer_1_weights[460][12] = 3;
        layer_1_weights[461][12] = 0;
        layer_1_weights[462][12] = 0;
        layer_1_weights[463][12] = -1;
        layer_1_weights[464][12] = -1;
        layer_1_weights[465][12] = 0;
        layer_1_weights[466][12] = -1;
        layer_1_weights[467][12] = -2;
        layer_1_weights[468][12] = -3;
        layer_1_weights[469][12] = -2;
        layer_1_weights[470][12] = -2;
        layer_1_weights[471][12] = -1;
        layer_1_weights[472][12] = -3;
        layer_1_weights[473][12] = -1;
        layer_1_weights[474][12] = -3;
        layer_1_weights[475][12] = -2;
        layer_1_weights[476][12] = 0;
        layer_1_weights[477][12] = -2;
        layer_1_weights[478][12] = -1;
        layer_1_weights[479][12] = 4;
        layer_1_weights[480][12] = -2;
        layer_1_weights[481][12] = -1;
        layer_1_weights[482][12] = 0;
        layer_1_weights[483][12] = -1;
        layer_1_weights[484][12] = -1;
        layer_1_weights[485][12] = 0;
        layer_1_weights[486][12] = 3;
        layer_1_weights[487][12] = 2;
        layer_1_weights[488][12] = 1;
        layer_1_weights[489][12] = 0;
        layer_1_weights[490][12] = -1;
        layer_1_weights[491][12] = 1;
        layer_1_weights[492][12] = 0;
        layer_1_weights[493][12] = 0;
        layer_1_weights[494][12] = 0;
        layer_1_weights[495][12] = -1;
        layer_1_weights[496][12] = 0;
        layer_1_weights[497][12] = 1;
        layer_1_weights[498][12] = -1;
        layer_1_weights[499][12] = -1;
        layer_1_weights[500][12] = -2;
        layer_1_weights[501][12] = -6;
        layer_1_weights[502][12] = -5;
        layer_1_weights[503][12] = -2;
        layer_1_weights[504][12] = -1;
        layer_1_weights[505][12] = 0;
        layer_1_weights[506][12] = -3;
        layer_1_weights[507][12] = -1;
        layer_1_weights[508][12] = -3;
        layer_1_weights[509][12] = 1;
        layer_1_weights[510][12] = -1;
        layer_1_weights[511][12] = -1;
        layer_1_weights[512][12] = 1;
        layer_1_weights[513][12] = 2;
        layer_1_weights[514][12] = 2;
        layer_1_weights[515][12] = 1;
        layer_1_weights[516][12] = 1;
        layer_1_weights[517][12] = 0;
        layer_1_weights[518][12] = -1;
        layer_1_weights[519][12] = 0;
        layer_1_weights[520][12] = 1;
        layer_1_weights[521][12] = 0;
        layer_1_weights[522][12] = -1;
        layer_1_weights[523][12] = -1;
        layer_1_weights[524][12] = -2;
        layer_1_weights[525][12] = -1;
        layer_1_weights[526][12] = -2;
        layer_1_weights[527][12] = -2;
        layer_1_weights[528][12] = -2;
        layer_1_weights[529][12] = 0;
        layer_1_weights[530][12] = -2;
        layer_1_weights[531][12] = -4;
        layer_1_weights[532][12] = -1;
        layer_1_weights[533][12] = -2;
        layer_1_weights[534][12] = -4;
        layer_1_weights[535][12] = -3;
        layer_1_weights[536][12] = -4;
        layer_1_weights[537][12] = 0;
        layer_1_weights[538][12] = 1;
        layer_1_weights[539][12] = -1;
        layer_1_weights[540][12] = 0;
        layer_1_weights[541][12] = 0;
        layer_1_weights[542][12] = 1;
        layer_1_weights[543][12] = 0;
        layer_1_weights[544][12] = 1;
        layer_1_weights[545][12] = 0;
        layer_1_weights[546][12] = 0;
        layer_1_weights[547][12] = -1;
        layer_1_weights[548][12] = -1;
        layer_1_weights[549][12] = -1;
        layer_1_weights[550][12] = 1;
        layer_1_weights[551][12] = -2;
        layer_1_weights[552][12] = -1;
        layer_1_weights[553][12] = -1;
        layer_1_weights[554][12] = 0;
        layer_1_weights[555][12] = -1;
        layer_1_weights[556][12] = 0;
        layer_1_weights[557][12] = 1;
        layer_1_weights[558][12] = 0;
        layer_1_weights[559][12] = -3;
        layer_1_weights[560][12] = 0;
        layer_1_weights[561][12] = -1;
        layer_1_weights[562][12] = -2;
        layer_1_weights[563][12] = -2;
        layer_1_weights[564][12] = -4;
        layer_1_weights[565][12] = -1;
        layer_1_weights[566][12] = -1;
        layer_1_weights[567][12] = -1;
        layer_1_weights[568][12] = 1;
        layer_1_weights[569][12] = 0;
        layer_1_weights[570][12] = 0;
        layer_1_weights[571][12] = 1;
        layer_1_weights[572][12] = 2;
        layer_1_weights[573][12] = 0;
        layer_1_weights[574][12] = 1;
        layer_1_weights[575][12] = -1;
        layer_1_weights[576][12] = -1;
        layer_1_weights[577][12] = -1;
        layer_1_weights[578][12] = -1;
        layer_1_weights[579][12] = 0;
        layer_1_weights[580][12] = 0;
        layer_1_weights[581][12] = 0;
        layer_1_weights[582][12] = -2;
        layer_1_weights[583][12] = 1;
        layer_1_weights[584][12] = -3;
        layer_1_weights[585][12] = 0;
        layer_1_weights[586][12] = -1;
        layer_1_weights[587][12] = 1;
        layer_1_weights[588][12] = 0;
        layer_1_weights[589][12] = -3;
        layer_1_weights[590][12] = -3;
        layer_1_weights[591][12] = -1;
        layer_1_weights[592][12] = -3;
        layer_1_weights[593][12] = -2;
        layer_1_weights[594][12] = -2;
        layer_1_weights[595][12] = -1;
        layer_1_weights[596][12] = 1;
        layer_1_weights[597][12] = 1;
        layer_1_weights[598][12] = 1;
        layer_1_weights[599][12] = 1;
        layer_1_weights[600][12] = 2;
        layer_1_weights[601][12] = 2;
        layer_1_weights[602][12] = 1;
        layer_1_weights[603][12] = 2;
        layer_1_weights[604][12] = 0;
        layer_1_weights[605][12] = 0;
        layer_1_weights[606][12] = 1;
        layer_1_weights[607][12] = 0;
        layer_1_weights[608][12] = 0;
        layer_1_weights[609][12] = 0;
        layer_1_weights[610][12] = 0;
        layer_1_weights[611][12] = -1;
        layer_1_weights[612][12] = -4;
        layer_1_weights[613][12] = 0;
        layer_1_weights[614][12] = -2;
        layer_1_weights[615][12] = -1;
        layer_1_weights[616][12] = 0;
        layer_1_weights[617][12] = 0;
        layer_1_weights[618][12] = -5;
        layer_1_weights[619][12] = 0;
        layer_1_weights[620][12] = 0;
        layer_1_weights[621][12] = -1;
        layer_1_weights[622][12] = -1;
        layer_1_weights[623][12] = -3;
        layer_1_weights[624][12] = -2;
        layer_1_weights[625][12] = -1;
        layer_1_weights[626][12] = 0;
        layer_1_weights[627][12] = 1;
        layer_1_weights[628][12] = 1;
        layer_1_weights[629][12] = 2;
        layer_1_weights[630][12] = 3;
        layer_1_weights[631][12] = 1;
        layer_1_weights[632][12] = 1;
        layer_1_weights[633][12] = 0;
        layer_1_weights[634][12] = -1;
        layer_1_weights[635][12] = 0;
        layer_1_weights[636][12] = 0;
        layer_1_weights[637][12] = -2;
        layer_1_weights[638][12] = -1;
        layer_1_weights[639][12] = 1;
        layer_1_weights[640][12] = 2;
        layer_1_weights[641][12] = 1;
        layer_1_weights[642][12] = 1;
        layer_1_weights[643][12] = -2;
        layer_1_weights[644][12] = -1;
        layer_1_weights[645][12] = 0;
        layer_1_weights[646][12] = -1;
        layer_1_weights[647][12] = 1;
        layer_1_weights[648][12] = -3;
        layer_1_weights[649][12] = -2;
        layer_1_weights[650][12] = -1;
        layer_1_weights[651][12] = -2;
        layer_1_weights[652][12] = -1;
        layer_1_weights[653][12] = -1;
        layer_1_weights[654][12] = -1;
        layer_1_weights[655][12] = 0;
        layer_1_weights[656][12] = 1;
        layer_1_weights[657][12] = 1;
        layer_1_weights[658][12] = 1;
        layer_1_weights[659][12] = 2;
        layer_1_weights[660][12] = 2;
        layer_1_weights[661][12] = 3;
        layer_1_weights[662][12] = 1;
        layer_1_weights[663][12] = 0;
        layer_1_weights[664][12] = 2;
        layer_1_weights[665][12] = -1;
        layer_1_weights[666][12] = -2;
        layer_1_weights[667][12] = 1;
        layer_1_weights[668][12] = 1;
        layer_1_weights[669][12] = 2;
        layer_1_weights[670][12] = -5;
        layer_1_weights[671][12] = 0;
        layer_1_weights[672][12] = 0;
        layer_1_weights[673][12] = 0;
        layer_1_weights[674][12] = -3;
        layer_1_weights[675][12] = 0;
        layer_1_weights[676][12] = 2;
        layer_1_weights[677][12] = 1;
        layer_1_weights[678][12] = -2;
        layer_1_weights[679][12] = -1;
        layer_1_weights[680][12] = 0;
        layer_1_weights[681][12] = 1;
        layer_1_weights[682][12] = 1;
        layer_1_weights[683][12] = -1;
        layer_1_weights[684][12] = 0;
        layer_1_weights[685][12] = 0;
        layer_1_weights[686][12] = 0;
        layer_1_weights[687][12] = 1;
        layer_1_weights[688][12] = 2;
        layer_1_weights[689][12] = 0;
        layer_1_weights[690][12] = 1;
        layer_1_weights[691][12] = 0;
        layer_1_weights[692][12] = 2;
        layer_1_weights[693][12] = -3;
        layer_1_weights[694][12] = -1;
        layer_1_weights[695][12] = -1;
        layer_1_weights[696][12] = -2;
        layer_1_weights[697][12] = -3;
        layer_1_weights[698][12] = -1;
        layer_1_weights[699][12] = -1;
        layer_1_weights[700][12] = -1;
        layer_1_weights[701][12] = 0;
        layer_1_weights[702][12] = 2;
        layer_1_weights[703][12] = 1;
        layer_1_weights[704][12] = -1;
        layer_1_weights[705][12] = -1;
        layer_1_weights[706][12] = -1;
        layer_1_weights[707][12] = 0;
        layer_1_weights[708][12] = 0;
        layer_1_weights[709][12] = 1;
        layer_1_weights[710][12] = 1;
        layer_1_weights[711][12] = 0;
        layer_1_weights[712][12] = 0;
        layer_1_weights[713][12] = -2;
        layer_1_weights[714][12] = -1;
        layer_1_weights[715][12] = 1;
        layer_1_weights[716][12] = 2;
        layer_1_weights[717][12] = 2;
        layer_1_weights[718][12] = 2;
        layer_1_weights[719][12] = 2;
        layer_1_weights[720][12] = 3;
        layer_1_weights[721][12] = 0;
        layer_1_weights[722][12] = 7;
        layer_1_weights[723][12] = 1;
        layer_1_weights[724][12] = 1;
        layer_1_weights[725][12] = 1;
        layer_1_weights[726][12] = -2;
        layer_1_weights[727][12] = 0;
        layer_1_weights[728][12] = 0;
        layer_1_weights[729][12] = 0;
        layer_1_weights[730][12] = 1;
        layer_1_weights[731][12] = 2;
        layer_1_weights[732][12] = 1;
        layer_1_weights[733][12] = -2;
        layer_1_weights[734][12] = 0;
        layer_1_weights[735][12] = 0;
        layer_1_weights[736][12] = 0;
        layer_1_weights[737][12] = 1;
        layer_1_weights[738][12] = -1;
        layer_1_weights[739][12] = 1;
        layer_1_weights[740][12] = 0;
        layer_1_weights[741][12] = -1;
        layer_1_weights[742][12] = 0;
        layer_1_weights[743][12] = 0;
        layer_1_weights[744][12] = -1;
        layer_1_weights[745][12] = 2;
        layer_1_weights[746][12] = 2;
        layer_1_weights[747][12] = -2;
        layer_1_weights[748][12] = -2;
        layer_1_weights[749][12] = -1;
        layer_1_weights[750][12] = 0;
        layer_1_weights[751][12] = 3;
        layer_1_weights[752][12] = 1;
        layer_1_weights[753][12] = 0;
        layer_1_weights[754][12] = 0;
        layer_1_weights[755][12] = 0;
        layer_1_weights[756][12] = 0;
        layer_1_weights[757][12] = 1;
        layer_1_weights[758][12] = 0;
        layer_1_weights[759][12] = 0;
        layer_1_weights[760][12] = -1;
        layer_1_weights[761][12] = -1;
        layer_1_weights[762][12] = 0;
        layer_1_weights[763][12] = -2;
        layer_1_weights[764][12] = -3;
        layer_1_weights[765][12] = 0;
        layer_1_weights[766][12] = 1;
        layer_1_weights[767][12] = 2;
        layer_1_weights[768][12] = 1;
        layer_1_weights[769][12] = 0;
        layer_1_weights[770][12] = 3;
        layer_1_weights[771][12] = 3;
        layer_1_weights[772][12] = 1;
        layer_1_weights[773][12] = 2;
        layer_1_weights[774][12] = 4;
        layer_1_weights[775][12] = 1;
        layer_1_weights[776][12] = -1;
        layer_1_weights[777][12] = -3;
        layer_1_weights[778][12] = -3;
        layer_1_weights[779][12] = 0;
        layer_1_weights[780][12] = 0;
        layer_1_weights[781][12] = 0;
        layer_1_weights[782][12] = 1;
        layer_1_weights[783][12] = 0;
        layer_1_weights[0][13] = 0;
        layer_1_weights[1][13] = 0;
        layer_1_weights[2][13] = -1;
        layer_1_weights[3][13] = 0;
        layer_1_weights[4][13] = -1;
        layer_1_weights[5][13] = 0;
        layer_1_weights[6][13] = 1;
        layer_1_weights[7][13] = 0;
        layer_1_weights[8][13] = 0;
        layer_1_weights[9][13] = 0;
        layer_1_weights[10][13] = 0;
        layer_1_weights[11][13] = -1;
        layer_1_weights[12][13] = 0;
        layer_1_weights[13][13] = 0;
        layer_1_weights[14][13] = 0;
        layer_1_weights[15][13] = 0;
        layer_1_weights[16][13] = 0;
        layer_1_weights[17][13] = 0;
        layer_1_weights[18][13] = 0;
        layer_1_weights[19][13] = 1;
        layer_1_weights[20][13] = -1;
        layer_1_weights[21][13] = 0;
        layer_1_weights[22][13] = 1;
        layer_1_weights[23][13] = 1;
        layer_1_weights[24][13] = 0;
        layer_1_weights[25][13] = 0;
        layer_1_weights[26][13] = 0;
        layer_1_weights[27][13] = 0;
        layer_1_weights[28][13] = 1;
        layer_1_weights[29][13] = 0;
        layer_1_weights[30][13] = 0;
        layer_1_weights[31][13] = 1;
        layer_1_weights[32][13] = 0;
        layer_1_weights[33][13] = 0;
        layer_1_weights[34][13] = 0;
        layer_1_weights[35][13] = 1;
        layer_1_weights[36][13] = 1;
        layer_1_weights[37][13] = 2;
        layer_1_weights[38][13] = 2;
        layer_1_weights[39][13] = 3;
        layer_1_weights[40][13] = 1;
        layer_1_weights[41][13] = 1;
        layer_1_weights[42][13] = -2;
        layer_1_weights[43][13] = 1;
        layer_1_weights[44][13] = 2;
        layer_1_weights[45][13] = 2;
        layer_1_weights[46][13] = 0;
        layer_1_weights[47][13] = 1;
        layer_1_weights[48][13] = 0;
        layer_1_weights[49][13] = 1;
        layer_1_weights[50][13] = 1;
        layer_1_weights[51][13] = 0;
        layer_1_weights[52][13] = 0;
        layer_1_weights[53][13] = 0;
        layer_1_weights[54][13] = 0;
        layer_1_weights[55][13] = 0;
        layer_1_weights[56][13] = 0;
        layer_1_weights[57][13] = 0;
        layer_1_weights[58][13] = 0;
        layer_1_weights[59][13] = 0;
        layer_1_weights[60][13] = 0;
        layer_1_weights[61][13] = 0;
        layer_1_weights[62][13] = 2;
        layer_1_weights[63][13] = 1;
        layer_1_weights[64][13] = 5;
        layer_1_weights[65][13] = 5;
        layer_1_weights[66][13] = 5;
        layer_1_weights[67][13] = 4;
        layer_1_weights[68][13] = 5;
        layer_1_weights[69][13] = 2;
        layer_1_weights[70][13] = 1;
        layer_1_weights[71][13] = 1;
        layer_1_weights[72][13] = -2;
        layer_1_weights[73][13] = -2;
        layer_1_weights[74][13] = -1;
        layer_1_weights[75][13] = 0;
        layer_1_weights[76][13] = 0;
        layer_1_weights[77][13] = 3;
        layer_1_weights[78][13] = 1;
        layer_1_weights[79][13] = 4;
        layer_1_weights[80][13] = 2;
        layer_1_weights[81][13] = 0;
        layer_1_weights[82][13] = 0;
        layer_1_weights[83][13] = 0;
        layer_1_weights[84][13] = 0;
        layer_1_weights[85][13] = -1;
        layer_1_weights[86][13] = 2;
        layer_1_weights[87][13] = 0;
        layer_1_weights[88][13] = 0;
        layer_1_weights[89][13] = 0;
        layer_1_weights[90][13] = 2;
        layer_1_weights[91][13] = 0;
        layer_1_weights[92][13] = -1;
        layer_1_weights[93][13] = 0;
        layer_1_weights[94][13] = -1;
        layer_1_weights[95][13] = -1;
        layer_1_weights[96][13] = 1;
        layer_1_weights[97][13] = 1;
        layer_1_weights[98][13] = -1;
        layer_1_weights[99][13] = -1;
        layer_1_weights[100][13] = -1;
        layer_1_weights[101][13] = -2;
        layer_1_weights[102][13] = -2;
        layer_1_weights[103][13] = 0;
        layer_1_weights[104][13] = 1;
        layer_1_weights[105][13] = -3;
        layer_1_weights[106][13] = 1;
        layer_1_weights[107][13] = 2;
        layer_1_weights[108][13] = 1;
        layer_1_weights[109][13] = -1;
        layer_1_weights[110][13] = -2;
        layer_1_weights[111][13] = 1;
        layer_1_weights[112][13] = 0;
        layer_1_weights[113][13] = 0;
        layer_1_weights[114][13] = 2;
        layer_1_weights[115][13] = 1;
        layer_1_weights[116][13] = 1;
        layer_1_weights[117][13] = 0;
        layer_1_weights[118][13] = 0;
        layer_1_weights[119][13] = -1;
        layer_1_weights[120][13] = 0;
        layer_1_weights[121][13] = -1;
        layer_1_weights[122][13] = -3;
        layer_1_weights[123][13] = -3;
        layer_1_weights[124][13] = 0;
        layer_1_weights[125][13] = 0;
        layer_1_weights[126][13] = -1;
        layer_1_weights[127][13] = -1;
        layer_1_weights[128][13] = -2;
        layer_1_weights[129][13] = 1;
        layer_1_weights[130][13] = 1;
        layer_1_weights[131][13] = 1;
        layer_1_weights[132][13] = 2;
        layer_1_weights[133][13] = -1;
        layer_1_weights[134][13] = 1;
        layer_1_weights[135][13] = -1;
        layer_1_weights[136][13] = -1;
        layer_1_weights[137][13] = 1;
        layer_1_weights[138][13] = 3;
        layer_1_weights[139][13] = 0;
        layer_1_weights[140][13] = 0;
        layer_1_weights[141][13] = -1;
        layer_1_weights[142][13] = 3;
        layer_1_weights[143][13] = -2;
        layer_1_weights[144][13] = 1;
        layer_1_weights[145][13] = -2;
        layer_1_weights[146][13] = -1;
        layer_1_weights[147][13] = -1;
        layer_1_weights[148][13] = 1;
        layer_1_weights[149][13] = -1;
        layer_1_weights[150][13] = 0;
        layer_1_weights[151][13] = 0;
        layer_1_weights[152][13] = -1;
        layer_1_weights[153][13] = -1;
        layer_1_weights[154][13] = -1;
        layer_1_weights[155][13] = 0;
        layer_1_weights[156][13] = 0;
        layer_1_weights[157][13] = 0;
        layer_1_weights[158][13] = -1;
        layer_1_weights[159][13] = 0;
        layer_1_weights[160][13] = 0;
        layer_1_weights[161][13] = 1;
        layer_1_weights[162][13] = 1;
        layer_1_weights[163][13] = 1;
        layer_1_weights[164][13] = 2;
        layer_1_weights[165][13] = 1;
        layer_1_weights[166][13] = 1;
        layer_1_weights[167][13] = -3;
        layer_1_weights[168][13] = 0;
        layer_1_weights[169][13] = 0;
        layer_1_weights[170][13] = -1;
        layer_1_weights[171][13] = 0;
        layer_1_weights[172][13] = 4;
        layer_1_weights[173][13] = -2;
        layer_1_weights[174][13] = 0;
        layer_1_weights[175][13] = 1;
        layer_1_weights[176][13] = 1;
        layer_1_weights[177][13] = 0;
        layer_1_weights[178][13] = -1;
        layer_1_weights[179][13] = -1;
        layer_1_weights[180][13] = -1;
        layer_1_weights[181][13] = 1;
        layer_1_weights[182][13] = 1;
        layer_1_weights[183][13] = 1;
        layer_1_weights[184][13] = 2;
        layer_1_weights[185][13] = 1;
        layer_1_weights[186][13] = 2;
        layer_1_weights[187][13] = 0;
        layer_1_weights[188][13] = 0;
        layer_1_weights[189][13] = 0;
        layer_1_weights[190][13] = -2;
        layer_1_weights[191][13] = 1;
        layer_1_weights[192][13] = -2;
        layer_1_weights[193][13] = 0;
        layer_1_weights[194][13] = 3;
        layer_1_weights[195][13] = 2;
        layer_1_weights[196][13] = 1;
        layer_1_weights[197][13] = 1;
        layer_1_weights[198][13] = -1;
        layer_1_weights[199][13] = 1;
        layer_1_weights[200][13] = 2;
        layer_1_weights[201][13] = 0;
        layer_1_weights[202][13] = 0;
        layer_1_weights[203][13] = 0;
        layer_1_weights[204][13] = -1;
        layer_1_weights[205][13] = 0;
        layer_1_weights[206][13] = -1;
        layer_1_weights[207][13] = 0;
        layer_1_weights[208][13] = 1;
        layer_1_weights[209][13] = 1;
        layer_1_weights[210][13] = 1;
        layer_1_weights[211][13] = 0;
        layer_1_weights[212][13] = 1;
        layer_1_weights[213][13] = 0;
        layer_1_weights[214][13] = 2;
        layer_1_weights[215][13] = 1;
        layer_1_weights[216][13] = 0;
        layer_1_weights[217][13] = 0;
        layer_1_weights[218][13] = 2;
        layer_1_weights[219][13] = 1;
        layer_1_weights[220][13] = -1;
        layer_1_weights[221][13] = -1;
        layer_1_weights[222][13] = -2;
        layer_1_weights[223][13] = 3;
        layer_1_weights[224][13] = -1;
        layer_1_weights[225][13] = 2;
        layer_1_weights[226][13] = 0;
        layer_1_weights[227][13] = 3;
        layer_1_weights[228][13] = 2;
        layer_1_weights[229][13] = 1;
        layer_1_weights[230][13] = 1;
        layer_1_weights[231][13] = 2;
        layer_1_weights[232][13] = 0;
        layer_1_weights[233][13] = 1;
        layer_1_weights[234][13] = 0;
        layer_1_weights[235][13] = 0;
        layer_1_weights[236][13] = -1;
        layer_1_weights[237][13] = 1;
        layer_1_weights[238][13] = 2;
        layer_1_weights[239][13] = 1;
        layer_1_weights[240][13] = 2;
        layer_1_weights[241][13] = 0;
        layer_1_weights[242][13] = -1;
        layer_1_weights[243][13] = 1;
        layer_1_weights[244][13] = 2;
        layer_1_weights[245][13] = 0;
        layer_1_weights[246][13] = 0;
        layer_1_weights[247][13] = 0;
        layer_1_weights[248][13] = -1;
        layer_1_weights[249][13] = -1;
        layer_1_weights[250][13] = 1;
        layer_1_weights[251][13] = 0;
        layer_1_weights[252][13] = 2;
        layer_1_weights[253][13] = 3;
        layer_1_weights[254][13] = 0;
        layer_1_weights[255][13] = 2;
        layer_1_weights[256][13] = 1;
        layer_1_weights[257][13] = 2;
        layer_1_weights[258][13] = -1;
        layer_1_weights[259][13] = 0;
        layer_1_weights[260][13] = -1;
        layer_1_weights[261][13] = 0;
        layer_1_weights[262][13] = 1;
        layer_1_weights[263][13] = 0;
        layer_1_weights[264][13] = 0;
        layer_1_weights[265][13] = 1;
        layer_1_weights[266][13] = 1;
        layer_1_weights[267][13] = 2;
        layer_1_weights[268][13] = 2;
        layer_1_weights[269][13] = 1;
        layer_1_weights[270][13] = 0;
        layer_1_weights[271][13] = 0;
        layer_1_weights[272][13] = 0;
        layer_1_weights[273][13] = 0;
        layer_1_weights[274][13] = 0;
        layer_1_weights[275][13] = 1;
        layer_1_weights[276][13] = -1;
        layer_1_weights[277][13] = -2;
        layer_1_weights[278][13] = 2;
        layer_1_weights[279][13] = 2;
        layer_1_weights[280][13] = 2;
        layer_1_weights[281][13] = 4;
        layer_1_weights[282][13] = -1;
        layer_1_weights[283][13] = 1;
        layer_1_weights[284][13] = -2;
        layer_1_weights[285][13] = 2;
        layer_1_weights[286][13] = -1;
        layer_1_weights[287][13] = 0;
        layer_1_weights[288][13] = 1;
        layer_1_weights[289][13] = 0;
        layer_1_weights[290][13] = 2;
        layer_1_weights[291][13] = 1;
        layer_1_weights[292][13] = 0;
        layer_1_weights[293][13] = 0;
        layer_1_weights[294][13] = 1;
        layer_1_weights[295][13] = 0;
        layer_1_weights[296][13] = 1;
        layer_1_weights[297][13] = 0;
        layer_1_weights[298][13] = 0;
        layer_1_weights[299][13] = 1;
        layer_1_weights[300][13] = 1;
        layer_1_weights[301][13] = 1;
        layer_1_weights[302][13] = 1;
        layer_1_weights[303][13] = 2;
        layer_1_weights[304][13] = 2;
        layer_1_weights[305][13] = 0;
        layer_1_weights[306][13] = -3;
        layer_1_weights[307][13] = 3;
        layer_1_weights[308][13] = 3;
        layer_1_weights[309][13] = 3;
        layer_1_weights[310][13] = 0;
        layer_1_weights[311][13] = 3;
        layer_1_weights[312][13] = 0;
        layer_1_weights[313][13] = 2;
        layer_1_weights[314][13] = 2;
        layer_1_weights[315][13] = 0;
        layer_1_weights[316][13] = 0;
        layer_1_weights[317][13] = 1;
        layer_1_weights[318][13] = 1;
        layer_1_weights[319][13] = 0;
        layer_1_weights[320][13] = 0;
        layer_1_weights[321][13] = -3;
        layer_1_weights[322][13] = -1;
        layer_1_weights[323][13] = 0;
        layer_1_weights[324][13] = 0;
        layer_1_weights[325][13] = 1;
        layer_1_weights[326][13] = -1;
        layer_1_weights[327][13] = 0;
        layer_1_weights[328][13] = 1;
        layer_1_weights[329][13] = 1;
        layer_1_weights[330][13] = -1;
        layer_1_weights[331][13] = 0;
        layer_1_weights[332][13] = -2;
        layer_1_weights[333][13] = -3;
        layer_1_weights[334][13] = -4;
        layer_1_weights[335][13] = -1;
        layer_1_weights[336][13] = 1;
        layer_1_weights[337][13] = 3;
        layer_1_weights[338][13] = 2;
        layer_1_weights[339][13] = 1;
        layer_1_weights[340][13] = 0;
        layer_1_weights[341][13] = 1;
        layer_1_weights[342][13] = 1;
        layer_1_weights[343][13] = 2;
        layer_1_weights[344][13] = 2;
        layer_1_weights[345][13] = 0;
        layer_1_weights[346][13] = -1;
        layer_1_weights[347][13] = -2;
        layer_1_weights[348][13] = -4;
        layer_1_weights[349][13] = -4;
        layer_1_weights[350][13] = -3;
        layer_1_weights[351][13] = -1;
        layer_1_weights[352][13] = -1;
        layer_1_weights[353][13] = 0;
        layer_1_weights[354][13] = 0;
        layer_1_weights[355][13] = 0;
        layer_1_weights[356][13] = 0;
        layer_1_weights[357][13] = 0;
        layer_1_weights[358][13] = 1;
        layer_1_weights[359][13] = -1;
        layer_1_weights[360][13] = -2;
        layer_1_weights[361][13] = -3;
        layer_1_weights[362][13] = -4;
        layer_1_weights[363][13] = 1;
        layer_1_weights[364][13] = 0;
        layer_1_weights[365][13] = 0;
        layer_1_weights[366][13] = 3;
        layer_1_weights[367][13] = 2;
        layer_1_weights[368][13] = -1;
        layer_1_weights[369][13] = 0;
        layer_1_weights[370][13] = -1;
        layer_1_weights[371][13] = -1;
        layer_1_weights[372][13] = -1;
        layer_1_weights[373][13] = -2;
        layer_1_weights[374][13] = -2;
        layer_1_weights[375][13] = -2;
        layer_1_weights[376][13] = -3;
        layer_1_weights[377][13] = -3;
        layer_1_weights[378][13] = -1;
        layer_1_weights[379][13] = -1;
        layer_1_weights[380][13] = 0;
        layer_1_weights[381][13] = 0;
        layer_1_weights[382][13] = 0;
        layer_1_weights[383][13] = 0;
        layer_1_weights[384][13] = -1;
        layer_1_weights[385][13] = 0;
        layer_1_weights[386][13] = 1;
        layer_1_weights[387][13] = -2;
        layer_1_weights[388][13] = -2;
        layer_1_weights[389][13] = -2;
        layer_1_weights[390][13] = -2;
        layer_1_weights[391][13] = 2;
        layer_1_weights[392][13] = -1;
        layer_1_weights[393][13] = -1;
        layer_1_weights[394][13] = 4;
        layer_1_weights[395][13] = 1;
        layer_1_weights[396][13] = -3;
        layer_1_weights[397][13] = -1;
        layer_1_weights[398][13] = -2;
        layer_1_weights[399][13] = -4;
        layer_1_weights[400][13] = -3;
        layer_1_weights[401][13] = -3;
        layer_1_weights[402][13] = -2;
        layer_1_weights[403][13] = -3;
        layer_1_weights[404][13] = -2;
        layer_1_weights[405][13] = 0;
        layer_1_weights[406][13] = 0;
        layer_1_weights[407][13] = -1;
        layer_1_weights[408][13] = -1;
        layer_1_weights[409][13] = -2;
        layer_1_weights[410][13] = 0;
        layer_1_weights[411][13] = 1;
        layer_1_weights[412][13] = -1;
        layer_1_weights[413][13] = 1;
        layer_1_weights[414][13] = -1;
        layer_1_weights[415][13] = -5;
        layer_1_weights[416][13] = -3;
        layer_1_weights[417][13] = -1;
        layer_1_weights[418][13] = 1;
        layer_1_weights[419][13] = 3;
        layer_1_weights[420][13] = -2;
        layer_1_weights[421][13] = 0;
        layer_1_weights[422][13] = -1;
        layer_1_weights[423][13] = -2;
        layer_1_weights[424][13] = -2;
        layer_1_weights[425][13] = -1;
        layer_1_weights[426][13] = -4;
        layer_1_weights[427][13] = -1;
        layer_1_weights[428][13] = -5;
        layer_1_weights[429][13] = -7;
        layer_1_weights[430][13] = -2;
        layer_1_weights[431][13] = -2;
        layer_1_weights[432][13] = 0;
        layer_1_weights[433][13] = 0;
        layer_1_weights[434][13] = 1;
        layer_1_weights[435][13] = -1;
        layer_1_weights[436][13] = -1;
        layer_1_weights[437][13] = 0;
        layer_1_weights[438][13] = 0;
        layer_1_weights[439][13] = -2;
        layer_1_weights[440][13] = -2;
        layer_1_weights[441][13] = -2;
        layer_1_weights[442][13] = -4;
        layer_1_weights[443][13] = -4;
        layer_1_weights[444][13] = -2;
        layer_1_weights[445][13] = -2;
        layer_1_weights[446][13] = 3;
        layer_1_weights[447][13] = 2;
        layer_1_weights[448][13] = 1;
        layer_1_weights[449][13] = 0;
        layer_1_weights[450][13] = 1;
        layer_1_weights[451][13] = -2;
        layer_1_weights[452][13] = -2;
        layer_1_weights[453][13] = -2;
        layer_1_weights[454][13] = -6;
        layer_1_weights[455][13] = -6;
        layer_1_weights[456][13] = -6;
        layer_1_weights[457][13] = -5;
        layer_1_weights[458][13] = -1;
        layer_1_weights[459][13] = 1;
        layer_1_weights[460][13] = 2;
        layer_1_weights[461][13] = 2;
        layer_1_weights[462][13] = 0;
        layer_1_weights[463][13] = -2;
        layer_1_weights[464][13] = -1;
        layer_1_weights[465][13] = -1;
        layer_1_weights[466][13] = -1;
        layer_1_weights[467][13] = -2;
        layer_1_weights[468][13] = -2;
        layer_1_weights[469][13] = -4;
        layer_1_weights[470][13] = -2;
        layer_1_weights[471][13] = -1;
        layer_1_weights[472][13] = 0;
        layer_1_weights[473][13] = 0;
        layer_1_weights[474][13] = 1;
        layer_1_weights[475][13] = 3;
        layer_1_weights[476][13] = 0;
        layer_1_weights[477][13] = 0;
        layer_1_weights[478][13] = 0;
        layer_1_weights[479][13] = -2;
        layer_1_weights[480][13] = -5;
        layer_1_weights[481][13] = -2;
        layer_1_weights[482][13] = -4;
        layer_1_weights[483][13] = -8;
        layer_1_weights[484][13] = -4;
        layer_1_weights[485][13] = -2;
        layer_1_weights[486][13] = 2;
        layer_1_weights[487][13] = 3;
        layer_1_weights[488][13] = 3;
        layer_1_weights[489][13] = 2;
        layer_1_weights[490][13] = -3;
        layer_1_weights[491][13] = -2;
        layer_1_weights[492][13] = -1;
        layer_1_weights[493][13] = -1;
        layer_1_weights[494][13] = -2;
        layer_1_weights[495][13] = -1;
        layer_1_weights[496][13] = -1;
        layer_1_weights[497][13] = -4;
        layer_1_weights[498][13] = -1;
        layer_1_weights[499][13] = -1;
        layer_1_weights[500][13] = 2;
        layer_1_weights[501][13] = 3;
        layer_1_weights[502][13] = 3;
        layer_1_weights[503][13] = 2;
        layer_1_weights[504][13] = 1;
        layer_1_weights[505][13] = 1;
        layer_1_weights[506][13] = -3;
        layer_1_weights[507][13] = -1;
        layer_1_weights[508][13] = -1;
        layer_1_weights[509][13] = -3;
        layer_1_weights[510][13] = -3;
        layer_1_weights[511][13] = -3;
        layer_1_weights[512][13] = -1;
        layer_1_weights[513][13] = 0;
        layer_1_weights[514][13] = 3;
        layer_1_weights[515][13] = 4;
        layer_1_weights[516][13] = 3;
        layer_1_weights[517][13] = 1;
        layer_1_weights[518][13] = -1;
        layer_1_weights[519][13] = -1;
        layer_1_weights[520][13] = -1;
        layer_1_weights[521][13] = -1;
        layer_1_weights[522][13] = 0;
        layer_1_weights[523][13] = -1;
        layer_1_weights[524][13] = -3;
        layer_1_weights[525][13] = -3;
        layer_1_weights[526][13] = 0;
        layer_1_weights[527][13] = 2;
        layer_1_weights[528][13] = 3;
        layer_1_weights[529][13] = 1;
        layer_1_weights[530][13] = 2;
        layer_1_weights[531][13] = 3;
        layer_1_weights[532][13] = 1;
        layer_1_weights[533][13] = 0;
        layer_1_weights[534][13] = -3;
        layer_1_weights[535][13] = -1;
        layer_1_weights[536][13] = 0;
        layer_1_weights[537][13] = -3;
        layer_1_weights[538][13] = -3;
        layer_1_weights[539][13] = -1;
        layer_1_weights[540][13] = 0;
        layer_1_weights[541][13] = 2;
        layer_1_weights[542][13] = 4;
        layer_1_weights[543][13] = 4;
        layer_1_weights[544][13] = 3;
        layer_1_weights[545][13] = 2;
        layer_1_weights[546][13] = 2;
        layer_1_weights[547][13] = -1;
        layer_1_weights[548][13] = 1;
        layer_1_weights[549][13] = 0;
        layer_1_weights[550][13] = -1;
        layer_1_weights[551][13] = -1;
        layer_1_weights[552][13] = 0;
        layer_1_weights[553][13] = -2;
        layer_1_weights[554][13] = 0;
        layer_1_weights[555][13] = 0;
        layer_1_weights[556][13] = 2;
        layer_1_weights[557][13] = 2;
        layer_1_weights[558][13] = 4;
        layer_1_weights[559][13] = 3;
        layer_1_weights[560][13] = -1;
        layer_1_weights[561][13] = 1;
        layer_1_weights[562][13] = 1;
        layer_1_weights[563][13] = 0;
        layer_1_weights[564][13] = -1;
        layer_1_weights[565][13] = -4;
        layer_1_weights[566][13] = -1;
        layer_1_weights[567][13] = -2;
        layer_1_weights[568][13] = -1;
        layer_1_weights[569][13] = 0;
        layer_1_weights[570][13] = 4;
        layer_1_weights[571][13] = 4;
        layer_1_weights[572][13] = 3;
        layer_1_weights[573][13] = 1;
        layer_1_weights[574][13] = 2;
        layer_1_weights[575][13] = 2;
        layer_1_weights[576][13] = 2;
        layer_1_weights[577][13] = 2;
        layer_1_weights[578][13] = 0;
        layer_1_weights[579][13] = 0;
        layer_1_weights[580][13] = 1;
        layer_1_weights[581][13] = 1;
        layer_1_weights[582][13] = 0;
        layer_1_weights[583][13] = -1;
        layer_1_weights[584][13] = 1;
        layer_1_weights[585][13] = 3;
        layer_1_weights[586][13] = 3;
        layer_1_weights[587][13] = 0;
        layer_1_weights[588][13] = 1;
        layer_1_weights[589][13] = 1;
        layer_1_weights[590][13] = 0;
        layer_1_weights[591][13] = -1;
        layer_1_weights[592][13] = -4;
        layer_1_weights[593][13] = -1;
        layer_1_weights[594][13] = -1;
        layer_1_weights[595][13] = -3;
        layer_1_weights[596][13] = -1;
        layer_1_weights[597][13] = -1;
        layer_1_weights[598][13] = 2;
        layer_1_weights[599][13] = 2;
        layer_1_weights[600][13] = 3;
        layer_1_weights[601][13] = 2;
        layer_1_weights[602][13] = 2;
        layer_1_weights[603][13] = 2;
        layer_1_weights[604][13] = 1;
        layer_1_weights[605][13] = 0;
        layer_1_weights[606][13] = 2;
        layer_1_weights[607][13] = 3;
        layer_1_weights[608][13] = 0;
        layer_1_weights[609][13] = -1;
        layer_1_weights[610][13] = 0;
        layer_1_weights[611][13] = 0;
        layer_1_weights[612][13] = 3;
        layer_1_weights[613][13] = 6;
        layer_1_weights[614][13] = 2;
        layer_1_weights[615][13] = 0;
        layer_1_weights[616][13] = 0;
        layer_1_weights[617][13] = 0;
        layer_1_weights[618][13] = 2;
        layer_1_weights[619][13] = -1;
        layer_1_weights[620][13] = 1;
        layer_1_weights[621][13] = -1;
        layer_1_weights[622][13] = 0;
        layer_1_weights[623][13] = 1;
        layer_1_weights[624][13] = 0;
        layer_1_weights[625][13] = 0;
        layer_1_weights[626][13] = -2;
        layer_1_weights[627][13] = 0;
        layer_1_weights[628][13] = 1;
        layer_1_weights[629][13] = 2;
        layer_1_weights[630][13] = 1;
        layer_1_weights[631][13] = 2;
        layer_1_weights[632][13] = 2;
        layer_1_weights[633][13] = 2;
        layer_1_weights[634][13] = 3;
        layer_1_weights[635][13] = 1;
        layer_1_weights[636][13] = 2;
        layer_1_weights[637][13] = 1;
        layer_1_weights[638][13] = 1;
        layer_1_weights[639][13] = 3;
        layer_1_weights[640][13] = 4;
        layer_1_weights[641][13] = 3;
        layer_1_weights[642][13] = 1;
        layer_1_weights[643][13] = -1;
        layer_1_weights[644][13] = 1;
        layer_1_weights[645][13] = 0;
        layer_1_weights[646][13] = -3;
        layer_1_weights[647][13] = -4;
        layer_1_weights[648][13] = 0;
        layer_1_weights[649][13] = 2;
        layer_1_weights[650][13] = 1;
        layer_1_weights[651][13] = 1;
        layer_1_weights[652][13] = 0;
        layer_1_weights[653][13] = 0;
        layer_1_weights[654][13] = -1;
        layer_1_weights[655][13] = 1;
        layer_1_weights[656][13] = 1;
        layer_1_weights[657][13] = 2;
        layer_1_weights[658][13] = 2;
        layer_1_weights[659][13] = 1;
        layer_1_weights[660][13] = 0;
        layer_1_weights[661][13] = -1;
        layer_1_weights[662][13] = 0;
        layer_1_weights[663][13] = 2;
        layer_1_weights[664][13] = 0;
        layer_1_weights[665][13] = 2;
        layer_1_weights[666][13] = 3;
        layer_1_weights[667][13] = 3;
        layer_1_weights[668][13] = 4;
        layer_1_weights[669][13] = 2;
        layer_1_weights[670][13] = 2;
        layer_1_weights[671][13] = 0;
        layer_1_weights[672][13] = 1;
        layer_1_weights[673][13] = 0;
        layer_1_weights[674][13] = 2;
        layer_1_weights[675][13] = 0;
        layer_1_weights[676][13] = -2;
        layer_1_weights[677][13] = -1;
        layer_1_weights[678][13] = -1;
        layer_1_weights[679][13] = -2;
        layer_1_weights[680][13] = -1;
        layer_1_weights[681][13] = -2;
        layer_1_weights[682][13] = -2;
        layer_1_weights[683][13] = 1;
        layer_1_weights[684][13] = 1;
        layer_1_weights[685][13] = 0;
        layer_1_weights[686][13] = 1;
        layer_1_weights[687][13] = 1;
        layer_1_weights[688][13] = 1;
        layer_1_weights[689][13] = 1;
        layer_1_weights[690][13] = 0;
        layer_1_weights[691][13] = 3;
        layer_1_weights[692][13] = 1;
        layer_1_weights[693][13] = 2;
        layer_1_weights[694][13] = 3;
        layer_1_weights[695][13] = 2;
        layer_1_weights[696][13] = 5;
        layer_1_weights[697][13] = 3;
        layer_1_weights[698][13] = 3;
        layer_1_weights[699][13] = 0;
        layer_1_weights[700][13] = -1;
        layer_1_weights[701][13] = 0;
        layer_1_weights[702][13] = -3;
        layer_1_weights[703][13] = 4;
        layer_1_weights[704][13] = -1;
        layer_1_weights[705][13] = -2;
        layer_1_weights[706][13] = 0;
        layer_1_weights[707][13] = -2;
        layer_1_weights[708][13] = 0;
        layer_1_weights[709][13] = -1;
        layer_1_weights[710][13] = -2;
        layer_1_weights[711][13] = -1;
        layer_1_weights[712][13] = 0;
        layer_1_weights[713][13] = -1;
        layer_1_weights[714][13] = 1;
        layer_1_weights[715][13] = 1;
        layer_1_weights[716][13] = 0;
        layer_1_weights[717][13] = 2;
        layer_1_weights[718][13] = 2;
        layer_1_weights[719][13] = 0;
        layer_1_weights[720][13] = 2;
        layer_1_weights[721][13] = 0;
        layer_1_weights[722][13] = 0;
        layer_1_weights[723][13] = -2;
        layer_1_weights[724][13] = 1;
        layer_1_weights[725][13] = 0;
        layer_1_weights[726][13] = 2;
        layer_1_weights[727][13] = 0;
        layer_1_weights[728][13] = 0;
        layer_1_weights[729][13] = 0;
        layer_1_weights[730][13] = 0;
        layer_1_weights[731][13] = 1;
        layer_1_weights[732][13] = -2;
        layer_1_weights[733][13] = -2;
        layer_1_weights[734][13] = 0;
        layer_1_weights[735][13] = 3;
        layer_1_weights[736][13] = 5;
        layer_1_weights[737][13] = 2;
        layer_1_weights[738][13] = 1;
        layer_1_weights[739][13] = 0;
        layer_1_weights[740][13] = 0;
        layer_1_weights[741][13] = 0;
        layer_1_weights[742][13] = -1;
        layer_1_weights[743][13] = -1;
        layer_1_weights[744][13] = 0;
        layer_1_weights[745][13] = -1;
        layer_1_weights[746][13] = 0;
        layer_1_weights[747][13] = 2;
        layer_1_weights[748][13] = 1;
        layer_1_weights[749][13] = 2;
        layer_1_weights[750][13] = 1;
        layer_1_weights[751][13] = 0;
        layer_1_weights[752][13] = 0;
        layer_1_weights[753][13] = 2;
        layer_1_weights[754][13] = 0;
        layer_1_weights[755][13] = 0;
        layer_1_weights[756][13] = 0;
        layer_1_weights[757][13] = 0;
        layer_1_weights[758][13] = 0;
        layer_1_weights[759][13] = 0;
        layer_1_weights[760][13] = 3;
        layer_1_weights[761][13] = 4;
        layer_1_weights[762][13] = 4;
        layer_1_weights[763][13] = 5;
        layer_1_weights[764][13] = 5;
        layer_1_weights[765][13] = 2;
        layer_1_weights[766][13] = 1;
        layer_1_weights[767][13] = 0;
        layer_1_weights[768][13] = 2;
        layer_1_weights[769][13] = 5;
        layer_1_weights[770][13] = 7;
        layer_1_weights[771][13] = 3;
        layer_1_weights[772][13] = 5;
        layer_1_weights[773][13] = 2;
        layer_1_weights[774][13] = 3;
        layer_1_weights[775][13] = 6;
        layer_1_weights[776][13] = 3;
        layer_1_weights[777][13] = 1;
        layer_1_weights[778][13] = 0;
        layer_1_weights[779][13] = 1;
        layer_1_weights[780][13] = 0;
        layer_1_weights[781][13] = 0;
        layer_1_weights[782][13] = 0;
        layer_1_weights[783][13] = 0;
        layer_1_weights[0][14] = -1;
        layer_1_weights[1][14] = 0;
        layer_1_weights[2][14] = 0;
        layer_1_weights[3][14] = 1;
        layer_1_weights[4][14] = 0;
        layer_1_weights[5][14] = 1;
        layer_1_weights[6][14] = 0;
        layer_1_weights[7][14] = 0;
        layer_1_weights[8][14] = 0;
        layer_1_weights[9][14] = 0;
        layer_1_weights[10][14] = 0;
        layer_1_weights[11][14] = 1;
        layer_1_weights[12][14] = 0;
        layer_1_weights[13][14] = 2;
        layer_1_weights[14][14] = 2;
        layer_1_weights[15][14] = 0;
        layer_1_weights[16][14] = 0;
        layer_1_weights[17][14] = -1;
        layer_1_weights[18][14] = -1;
        layer_1_weights[19][14] = 0;
        layer_1_weights[20][14] = 0;
        layer_1_weights[21][14] = 0;
        layer_1_weights[22][14] = 0;
        layer_1_weights[23][14] = 0;
        layer_1_weights[24][14] = -1;
        layer_1_weights[25][14] = 1;
        layer_1_weights[26][14] = 0;
        layer_1_weights[27][14] = 1;
        layer_1_weights[28][14] = 0;
        layer_1_weights[29][14] = 0;
        layer_1_weights[30][14] = 0;
        layer_1_weights[31][14] = 0;
        layer_1_weights[32][14] = 0;
        layer_1_weights[33][14] = 1;
        layer_1_weights[34][14] = 0;
        layer_1_weights[35][14] = -2;
        layer_1_weights[36][14] = -2;
        layer_1_weights[37][14] = -2;
        layer_1_weights[38][14] = -1;
        layer_1_weights[39][14] = -3;
        layer_1_weights[40][14] = -4;
        layer_1_weights[41][14] = -1;
        layer_1_weights[42][14] = -3;
        layer_1_weights[43][14] = 4;
        layer_1_weights[44][14] = 4;
        layer_1_weights[45][14] = 3;
        layer_1_weights[46][14] = 2;
        layer_1_weights[47][14] = 3;
        layer_1_weights[48][14] = 3;
        layer_1_weights[49][14] = 1;
        layer_1_weights[50][14] = 3;
        layer_1_weights[51][14] = 1;
        layer_1_weights[52][14] = 1;
        layer_1_weights[53][14] = -1;
        layer_1_weights[54][14] = 0;
        layer_1_weights[55][14] = 0;
        layer_1_weights[56][14] = 0;
        layer_1_weights[57][14] = 0;
        layer_1_weights[58][14] = 2;
        layer_1_weights[59][14] = 0;
        layer_1_weights[60][14] = 0;
        layer_1_weights[61][14] = 1;
        layer_1_weights[62][14] = -4;
        layer_1_weights[63][14] = -1;
        layer_1_weights[64][14] = 3;
        layer_1_weights[65][14] = 5;
        layer_1_weights[66][14] = 3;
        layer_1_weights[67][14] = -1;
        layer_1_weights[68][14] = 1;
        layer_1_weights[69][14] = -2;
        layer_1_weights[70][14] = -3;
        layer_1_weights[71][14] = -2;
        layer_1_weights[72][14] = -1;
        layer_1_weights[73][14] = -2;
        layer_1_weights[74][14] = -1;
        layer_1_weights[75][14] = -3;
        layer_1_weights[76][14] = -1;
        layer_1_weights[77][14] = 2;
        layer_1_weights[78][14] = -1;
        layer_1_weights[79][14] = 1;
        layer_1_weights[80][14] = 5;
        layer_1_weights[81][14] = 2;
        layer_1_weights[82][14] = 0;
        layer_1_weights[83][14] = 1;
        layer_1_weights[84][14] = 0;
        layer_1_weights[85][14] = 0;
        layer_1_weights[86][14] = -3;
        layer_1_weights[87][14] = 3;
        layer_1_weights[88][14] = -3;
        layer_1_weights[89][14] = -1;
        layer_1_weights[90][14] = 2;
        layer_1_weights[91][14] = 0;
        layer_1_weights[92][14] = 1;
        layer_1_weights[93][14] = 1;
        layer_1_weights[94][14] = 3;
        layer_1_weights[95][14] = 2;
        layer_1_weights[96][14] = 1;
        layer_1_weights[97][14] = 1;
        layer_1_weights[98][14] = 3;
        layer_1_weights[99][14] = -1;
        layer_1_weights[100][14] = 0;
        layer_1_weights[101][14] = 0;
        layer_1_weights[102][14] = 0;
        layer_1_weights[103][14] = 0;
        layer_1_weights[104][14] = -2;
        layer_1_weights[105][14] = -2;
        layer_1_weights[106][14] = 0;
        layer_1_weights[107][14] = 2;
        layer_1_weights[108][14] = -1;
        layer_1_weights[109][14] = 2;
        layer_1_weights[110][14] = 0;
        layer_1_weights[111][14] = 0;
        layer_1_weights[112][14] = 0;
        layer_1_weights[113][14] = -1;
        layer_1_weights[114][14] = -3;
        layer_1_weights[115][14] = -4;
        layer_1_weights[116][14] = 0;
        layer_1_weights[117][14] = 0;
        layer_1_weights[118][14] = 1;
        layer_1_weights[119][14] = 0;
        layer_1_weights[120][14] = 2;
        layer_1_weights[121][14] = 3;
        layer_1_weights[122][14] = 1;
        layer_1_weights[123][14] = 0;
        layer_1_weights[124][14] = 2;
        layer_1_weights[125][14] = 2;
        layer_1_weights[126][14] = 2;
        layer_1_weights[127][14] = 2;
        layer_1_weights[128][14] = 2;
        layer_1_weights[129][14] = 3;
        layer_1_weights[130][14] = 1;
        layer_1_weights[131][14] = 0;
        layer_1_weights[132][14] = 0;
        layer_1_weights[133][14] = -1;
        layer_1_weights[134][14] = -1;
        layer_1_weights[135][14] = -2;
        layer_1_weights[136][14] = -2;
        layer_1_weights[137][14] = 0;
        layer_1_weights[138][14] = 2;
        layer_1_weights[139][14] = 3;
        layer_1_weights[140][14] = 0;
        layer_1_weights[141][14] = 1;
        layer_1_weights[142][14] = 4;
        layer_1_weights[143][14] = -4;
        layer_1_weights[144][14] = 1;
        layer_1_weights[145][14] = -2;
        layer_1_weights[146][14] = 1;
        layer_1_weights[147][14] = -3;
        layer_1_weights[148][14] = 0;
        layer_1_weights[149][14] = 1;
        layer_1_weights[150][14] = 1;
        layer_1_weights[151][14] = 2;
        layer_1_weights[152][14] = 1;
        layer_1_weights[153][14] = 1;
        layer_1_weights[154][14] = 1;
        layer_1_weights[155][14] = 2;
        layer_1_weights[156][14] = 3;
        layer_1_weights[157][14] = 2;
        layer_1_weights[158][14] = 2;
        layer_1_weights[159][14] = 1;
        layer_1_weights[160][14] = 1;
        layer_1_weights[161][14] = 2;
        layer_1_weights[162][14] = 1;
        layer_1_weights[163][14] = -2;
        layer_1_weights[164][14] = -3;
        layer_1_weights[165][14] = 0;
        layer_1_weights[166][14] = 0;
        layer_1_weights[167][14] = 0;
        layer_1_weights[168][14] = -1;
        layer_1_weights[169][14] = -1;
        layer_1_weights[170][14] = -3;
        layer_1_weights[171][14] = -2;
        layer_1_weights[172][14] = 1;
        layer_1_weights[173][14] = -2;
        layer_1_weights[174][14] = 0;
        layer_1_weights[175][14] = 0;
        layer_1_weights[176][14] = 0;
        layer_1_weights[177][14] = -1;
        layer_1_weights[178][14] = 0;
        layer_1_weights[179][14] = 1;
        layer_1_weights[180][14] = 0;
        layer_1_weights[181][14] = 0;
        layer_1_weights[182][14] = 0;
        layer_1_weights[183][14] = 0;
        layer_1_weights[184][14] = 1;
        layer_1_weights[185][14] = 0;
        layer_1_weights[186][14] = 1;
        layer_1_weights[187][14] = 1;
        layer_1_weights[188][14] = 1;
        layer_1_weights[189][14] = 1;
        layer_1_weights[190][14] = 0;
        layer_1_weights[191][14] = -1;
        layer_1_weights[192][14] = -4;
        layer_1_weights[193][14] = 1;
        layer_1_weights[194][14] = -2;
        layer_1_weights[195][14] = 1;
        layer_1_weights[196][14] = -1;
        layer_1_weights[197][14] = -3;
        layer_1_weights[198][14] = -2;
        layer_1_weights[199][14] = -1;
        layer_1_weights[200][14] = 2;
        layer_1_weights[201][14] = 0;
        layer_1_weights[202][14] = -1;
        layer_1_weights[203][14] = 1;
        layer_1_weights[204][14] = 0;
        layer_1_weights[205][14] = 1;
        layer_1_weights[206][14] = 0;
        layer_1_weights[207][14] = 0;
        layer_1_weights[208][14] = -1;
        layer_1_weights[209][14] = 0;
        layer_1_weights[210][14] = -1;
        layer_1_weights[211][14] = 0;
        layer_1_weights[212][14] = 0;
        layer_1_weights[213][14] = 1;
        layer_1_weights[214][14] = 0;
        layer_1_weights[215][14] = 1;
        layer_1_weights[216][14] = -1;
        layer_1_weights[217][14] = 0;
        layer_1_weights[218][14] = 1;
        layer_1_weights[219][14] = -1;
        layer_1_weights[220][14] = -1;
        layer_1_weights[221][14] = 0;
        layer_1_weights[222][14] = -2;
        layer_1_weights[223][14] = 2;
        layer_1_weights[224][14] = 2;
        layer_1_weights[225][14] = 1;
        layer_1_weights[226][14] = 0;
        layer_1_weights[227][14] = 0;
        layer_1_weights[228][14] = -1;
        layer_1_weights[229][14] = 0;
        layer_1_weights[230][14] = 2;
        layer_1_weights[231][14] = 1;
        layer_1_weights[232][14] = 0;
        layer_1_weights[233][14] = 1;
        layer_1_weights[234][14] = 1;
        layer_1_weights[235][14] = 0;
        layer_1_weights[236][14] = 0;
        layer_1_weights[237][14] = 0;
        layer_1_weights[238][14] = 1;
        layer_1_weights[239][14] = -1;
        layer_1_weights[240][14] = 0;
        layer_1_weights[241][14] = 1;
        layer_1_weights[242][14] = 0;
        layer_1_weights[243][14] = 1;
        layer_1_weights[244][14] = 1;
        layer_1_weights[245][14] = 0;
        layer_1_weights[246][14] = 1;
        layer_1_weights[247][14] = -1;
        layer_1_weights[248][14] = -2;
        layer_1_weights[249][14] = -1;
        layer_1_weights[250][14] = 1;
        layer_1_weights[251][14] = -1;
        layer_1_weights[252][14] = -1;
        layer_1_weights[253][14] = -3;
        layer_1_weights[254][14] = -1;
        layer_1_weights[255][14] = 0;
        layer_1_weights[256][14] = 1;
        layer_1_weights[257][14] = 1;
        layer_1_weights[258][14] = -1;
        layer_1_weights[259][14] = -1;
        layer_1_weights[260][14] = 0;
        layer_1_weights[261][14] = 1;
        layer_1_weights[262][14] = 0;
        layer_1_weights[263][14] = 0;
        layer_1_weights[264][14] = -1;
        layer_1_weights[265][14] = 0;
        layer_1_weights[266][14] = -2;
        layer_1_weights[267][14] = 1;
        layer_1_weights[268][14] = 0;
        layer_1_weights[269][14] = 0;
        layer_1_weights[270][14] = 0;
        layer_1_weights[271][14] = 1;
        layer_1_weights[272][14] = 0;
        layer_1_weights[273][14] = 1;
        layer_1_weights[274][14] = -1;
        layer_1_weights[275][14] = -2;
        layer_1_weights[276][14] = -2;
        layer_1_weights[277][14] = -3;
        layer_1_weights[278][14] = -1;
        layer_1_weights[279][14] = -2;
        layer_1_weights[280][14] = 0;
        layer_1_weights[281][14] = -2;
        layer_1_weights[282][14] = -1;
        layer_1_weights[283][14] = 0;
        layer_1_weights[284][14] = 0;
        layer_1_weights[285][14] = 2;
        layer_1_weights[286][14] = 0;
        layer_1_weights[287][14] = 1;
        layer_1_weights[288][14] = 1;
        layer_1_weights[289][14] = 0;
        layer_1_weights[290][14] = -1;
        layer_1_weights[291][14] = 0;
        layer_1_weights[292][14] = 0;
        layer_1_weights[293][14] = -1;
        layer_1_weights[294][14] = 0;
        layer_1_weights[295][14] = -2;
        layer_1_weights[296][14] = -2;
        layer_1_weights[297][14] = -1;
        layer_1_weights[298][14] = 1;
        layer_1_weights[299][14] = 1;
        layer_1_weights[300][14] = 2;
        layer_1_weights[301][14] = 1;
        layer_1_weights[302][14] = -2;
        layer_1_weights[303][14] = 1;
        layer_1_weights[304][14] = -2;
        layer_1_weights[305][14] = -4;
        layer_1_weights[306][14] = -2;
        layer_1_weights[307][14] = -2;
        layer_1_weights[308][14] = -2;
        layer_1_weights[309][14] = 1;
        layer_1_weights[310][14] = 0;
        layer_1_weights[311][14] = 0;
        layer_1_weights[312][14] = -1;
        layer_1_weights[313][14] = 3;
        layer_1_weights[314][14] = 1;
        layer_1_weights[315][14] = 0;
        layer_1_weights[316][14] = 0;
        layer_1_weights[317][14] = 0;
        layer_1_weights[318][14] = -1;
        layer_1_weights[319][14] = -1;
        layer_1_weights[320][14] = 0;
        layer_1_weights[321][14] = -3;
        layer_1_weights[322][14] = -3;
        layer_1_weights[323][14] = -3;
        layer_1_weights[324][14] = -3;
        layer_1_weights[325][14] = -1;
        layer_1_weights[326][14] = -1;
        layer_1_weights[327][14] = 1;
        layer_1_weights[328][14] = 1;
        layer_1_weights[329][14] = 0;
        layer_1_weights[330][14] = 1;
        layer_1_weights[331][14] = 0;
        layer_1_weights[332][14] = 1;
        layer_1_weights[333][14] = -1;
        layer_1_weights[334][14] = 2;
        layer_1_weights[335][14] = 1;
        layer_1_weights[336][14] = -2;
        layer_1_weights[337][14] = -1;
        layer_1_weights[338][14] = -1;
        layer_1_weights[339][14] = 0;
        layer_1_weights[340][14] = 2;
        layer_1_weights[341][14] = 1;
        layer_1_weights[342][14] = -1;
        layer_1_weights[343][14] = 0;
        layer_1_weights[344][14] = 0;
        layer_1_weights[345][14] = 1;
        layer_1_weights[346][14] = -1;
        layer_1_weights[347][14] = -1;
        layer_1_weights[348][14] = 0;
        layer_1_weights[349][14] = 0;
        layer_1_weights[350][14] = -3;
        layer_1_weights[351][14] = -3;
        layer_1_weights[352][14] = -1;
        layer_1_weights[353][14] = -2;
        layer_1_weights[354][14] = 0;
        layer_1_weights[355][14] = 1;
        layer_1_weights[356][14] = 1;
        layer_1_weights[357][14] = 2;
        layer_1_weights[358][14] = 0;
        layer_1_weights[359][14] = 0;
        layer_1_weights[360][14] = 3;
        layer_1_weights[361][14] = 0;
        layer_1_weights[362][14] = -1;
        layer_1_weights[363][14] = -2;
        layer_1_weights[364][14] = 0;
        layer_1_weights[365][14] = 2;
        layer_1_weights[366][14] = 1;
        layer_1_weights[367][14] = -1;
        layer_1_weights[368][14] = 0;
        layer_1_weights[369][14] = 1;
        layer_1_weights[370][14] = 2;
        layer_1_weights[371][14] = 1;
        layer_1_weights[372][14] = -1;
        layer_1_weights[373][14] = -2;
        layer_1_weights[374][14] = 0;
        layer_1_weights[375][14] = 1;
        layer_1_weights[376][14] = 2;
        layer_1_weights[377][14] = 1;
        layer_1_weights[378][14] = 0;
        layer_1_weights[379][14] = 0;
        layer_1_weights[380][14] = 0;
        layer_1_weights[381][14] = 0;
        layer_1_weights[382][14] = 0;
        layer_1_weights[383][14] = 1;
        layer_1_weights[384][14] = 1;
        layer_1_weights[385][14] = 1;
        layer_1_weights[386][14] = 3;
        layer_1_weights[387][14] = 3;
        layer_1_weights[388][14] = 6;
        layer_1_weights[389][14] = 1;
        layer_1_weights[390][14] = 1;
        layer_1_weights[391][14] = 3;
        layer_1_weights[392][14] = -2;
        layer_1_weights[393][14] = -1;
        layer_1_weights[394][14] = -5;
        layer_1_weights[395][14] = -2;
        layer_1_weights[396][14] = 0;
        layer_1_weights[397][14] = 0;
        layer_1_weights[398][14] = 0;
        layer_1_weights[399][14] = 0;
        layer_1_weights[400][14] = 0;
        layer_1_weights[401][14] = 1;
        layer_1_weights[402][14] = 2;
        layer_1_weights[403][14] = 1;
        layer_1_weights[404][14] = 3;
        layer_1_weights[405][14] = 3;
        layer_1_weights[406][14] = 2;
        layer_1_weights[407][14] = 1;
        layer_1_weights[408][14] = 0;
        layer_1_weights[409][14] = 0;
        layer_1_weights[410][14] = 0;
        layer_1_weights[411][14] = 0;
        layer_1_weights[412][14] = -1;
        layer_1_weights[413][14] = -1;
        layer_1_weights[414][14] = -1;
        layer_1_weights[415][14] = 0;
        layer_1_weights[416][14] = 1;
        layer_1_weights[417][14] = 5;
        layer_1_weights[418][14] = 3;
        layer_1_weights[419][14] = 2;
        layer_1_weights[420][14] = -2;
        layer_1_weights[421][14] = -1;
        layer_1_weights[422][14] = 0;
        layer_1_weights[423][14] = 0;
        layer_1_weights[424][14] = 1;
        layer_1_weights[425][14] = 1;
        layer_1_weights[426][14] = 1;
        layer_1_weights[427][14] = 0;
        layer_1_weights[428][14] = 1;
        layer_1_weights[429][14] = 0;
        layer_1_weights[430][14] = 2;
        layer_1_weights[431][14] = 2;
        layer_1_weights[432][14] = 2;
        layer_1_weights[433][14] = 2;
        layer_1_weights[434][14] = 1;
        layer_1_weights[435][14] = 1;
        layer_1_weights[436][14] = 1;
        layer_1_weights[437][14] = 0;
        layer_1_weights[438][14] = 1;
        layer_1_weights[439][14] = 1;
        layer_1_weights[440][14] = -1;
        layer_1_weights[441][14] = -1;
        layer_1_weights[442][14] = -1;
        layer_1_weights[443][14] = -1;
        layer_1_weights[444][14] = 3;
        layer_1_weights[445][14] = 2;
        layer_1_weights[446][14] = 3;
        layer_1_weights[447][14] = 4;
        layer_1_weights[448][14] = -1;
        layer_1_weights[449][14] = -1;
        layer_1_weights[450][14] = 2;
        layer_1_weights[451][14] = 1;
        layer_1_weights[452][14] = 0;
        layer_1_weights[453][14] = 0;
        layer_1_weights[454][14] = 0;
        layer_1_weights[455][14] = 1;
        layer_1_weights[456][14] = 1;
        layer_1_weights[457][14] = 3;
        layer_1_weights[458][14] = 3;
        layer_1_weights[459][14] = 2;
        layer_1_weights[460][14] = 1;
        layer_1_weights[461][14] = 2;
        layer_1_weights[462][14] = 1;
        layer_1_weights[463][14] = 1;
        layer_1_weights[464][14] = 2;
        layer_1_weights[465][14] = 1;
        layer_1_weights[466][14] = 0;
        layer_1_weights[467][14] = 1;
        layer_1_weights[468][14] = -1;
        layer_1_weights[469][14] = -1;
        layer_1_weights[470][14] = 1;
        layer_1_weights[471][14] = 1;
        layer_1_weights[472][14] = 1;
        layer_1_weights[473][14] = 5;
        layer_1_weights[474][14] = 6;
        layer_1_weights[475][14] = 4;
        layer_1_weights[476][14] = 0;
        layer_1_weights[477][14] = -2;
        layer_1_weights[478][14] = 1;
        layer_1_weights[479][14] = -2;
        layer_1_weights[480][14] = 0;
        layer_1_weights[481][14] = 1;
        layer_1_weights[482][14] = 1;
        layer_1_weights[483][14] = 0;
        layer_1_weights[484][14] = 1;
        layer_1_weights[485][14] = 3;
        layer_1_weights[486][14] = 2;
        layer_1_weights[487][14] = 2;
        layer_1_weights[488][14] = 2;
        layer_1_weights[489][14] = 1;
        layer_1_weights[490][14] = 0;
        layer_1_weights[491][14] = 1;
        layer_1_weights[492][14] = 2;
        layer_1_weights[493][14] = 1;
        layer_1_weights[494][14] = 0;
        layer_1_weights[495][14] = -1;
        layer_1_weights[496][14] = 0;
        layer_1_weights[497][14] = 1;
        layer_1_weights[498][14] = 1;
        layer_1_weights[499][14] = 0;
        layer_1_weights[500][14] = -2;
        layer_1_weights[501][14] = 3;
        layer_1_weights[502][14] = 1;
        layer_1_weights[503][14] = 5;
        layer_1_weights[504][14] = 1;
        layer_1_weights[505][14] = -1;
        layer_1_weights[506][14] = -1;
        layer_1_weights[507][14] = -1;
        layer_1_weights[508][14] = 0;
        layer_1_weights[509][14] = -1;
        layer_1_weights[510][14] = 0;
        layer_1_weights[511][14] = 0;
        layer_1_weights[512][14] = 3;
        layer_1_weights[513][14] = 0;
        layer_1_weights[514][14] = 0;
        layer_1_weights[515][14] = -1;
        layer_1_weights[516][14] = 0;
        layer_1_weights[517][14] = 0;
        layer_1_weights[518][14] = 0;
        layer_1_weights[519][14] = 0;
        layer_1_weights[520][14] = -1;
        layer_1_weights[521][14] = 0;
        layer_1_weights[522][14] = -1;
        layer_1_weights[523][14] = 0;
        layer_1_weights[524][14] = 1;
        layer_1_weights[525][14] = 0;
        layer_1_weights[526][14] = 0;
        layer_1_weights[527][14] = 2;
        layer_1_weights[528][14] = 2;
        layer_1_weights[529][14] = 2;
        layer_1_weights[530][14] = -1;
        layer_1_weights[531][14] = 2;
        layer_1_weights[532][14] = 0;
        layer_1_weights[533][14] = 0;
        layer_1_weights[534][14] = -3;
        layer_1_weights[535][14] = -1;
        layer_1_weights[536][14] = 0;
        layer_1_weights[537][14] = 1;
        layer_1_weights[538][14] = 1;
        layer_1_weights[539][14] = 3;
        layer_1_weights[540][14] = 0;
        layer_1_weights[541][14] = 0;
        layer_1_weights[542][14] = 1;
        layer_1_weights[543][14] = -1;
        layer_1_weights[544][14] = -1;
        layer_1_weights[545][14] = 0;
        layer_1_weights[546][14] = 1;
        layer_1_weights[547][14] = 1;
        layer_1_weights[548][14] = 0;
        layer_1_weights[549][14] = 2;
        layer_1_weights[550][14] = 0;
        layer_1_weights[551][14] = 0;
        layer_1_weights[552][14] = 1;
        layer_1_weights[553][14] = 1;
        layer_1_weights[554][14] = 2;
        layer_1_weights[555][14] = 3;
        layer_1_weights[556][14] = 0;
        layer_1_weights[557][14] = -3;
        layer_1_weights[558][14] = 5;
        layer_1_weights[559][14] = 0;
        layer_1_weights[560][14] = 1;
        layer_1_weights[561][14] = 1;
        layer_1_weights[562][14] = 3;
        layer_1_weights[563][14] = 1;
        layer_1_weights[564][14] = 1;
        layer_1_weights[565][14] = -1;
        layer_1_weights[566][14] = 3;
        layer_1_weights[567][14] = 2;
        layer_1_weights[568][14] = 0;
        layer_1_weights[569][14] = 0;
        layer_1_weights[570][14] = 1;
        layer_1_weights[571][14] = 0;
        layer_1_weights[572][14] = 1;
        layer_1_weights[573][14] = -1;
        layer_1_weights[574][14] = 0;
        layer_1_weights[575][14] = 1;
        layer_1_weights[576][14] = 0;
        layer_1_weights[577][14] = 0;
        layer_1_weights[578][14] = 1;
        layer_1_weights[579][14] = 1;
        layer_1_weights[580][14] = 0;
        layer_1_weights[581][14] = 3;
        layer_1_weights[582][14] = 2;
        layer_1_weights[583][14] = 2;
        layer_1_weights[584][14] = 0;
        layer_1_weights[585][14] = -1;
        layer_1_weights[586][14] = 5;
        layer_1_weights[587][14] = -3;
        layer_1_weights[588][14] = 0;
        layer_1_weights[589][14] = 1;
        layer_1_weights[590][14] = 1;
        layer_1_weights[591][14] = 1;
        layer_1_weights[592][14] = 1;
        layer_1_weights[593][14] = 2;
        layer_1_weights[594][14] = 2;
        layer_1_weights[595][14] = 2;
        layer_1_weights[596][14] = 1;
        layer_1_weights[597][14] = 2;
        layer_1_weights[598][14] = 1;
        layer_1_weights[599][14] = 1;
        layer_1_weights[600][14] = 0;
        layer_1_weights[601][14] = 1;
        layer_1_weights[602][14] = -1;
        layer_1_weights[603][14] = 1;
        layer_1_weights[604][14] = 0;
        layer_1_weights[605][14] = -1;
        layer_1_weights[606][14] = 0;
        layer_1_weights[607][14] = 0;
        layer_1_weights[608][14] = 0;
        layer_1_weights[609][14] = 0;
        layer_1_weights[610][14] = 2;
        layer_1_weights[611][14] = 1;
        layer_1_weights[612][14] = -1;
        layer_1_weights[613][14] = -2;
        layer_1_weights[614][14] = 5;
        layer_1_weights[615][14] = 0;
        layer_1_weights[616][14] = 0;
        layer_1_weights[617][14] = -1;
        layer_1_weights[618][14] = 1;
        layer_1_weights[619][14] = 2;
        layer_1_weights[620][14] = 2;
        layer_1_weights[621][14] = 3;
        layer_1_weights[622][14] = 1;
        layer_1_weights[623][14] = 2;
        layer_1_weights[624][14] = 3;
        layer_1_weights[625][14] = 1;
        layer_1_weights[626][14] = 2;
        layer_1_weights[627][14] = 2;
        layer_1_weights[628][14] = 2;
        layer_1_weights[629][14] = 2;
        layer_1_weights[630][14] = 0;
        layer_1_weights[631][14] = -1;
        layer_1_weights[632][14] = -1;
        layer_1_weights[633][14] = 0;
        layer_1_weights[634][14] = 0;
        layer_1_weights[635][14] = 0;
        layer_1_weights[636][14] = 1;
        layer_1_weights[637][14] = 1;
        layer_1_weights[638][14] = 3;
        layer_1_weights[639][14] = 0;
        layer_1_weights[640][14] = -1;
        layer_1_weights[641][14] = -2;
        layer_1_weights[642][14] = -2;
        layer_1_weights[643][14] = -1;
        layer_1_weights[644][14] = 1;
        layer_1_weights[645][14] = 0;
        layer_1_weights[646][14] = 1;
        layer_1_weights[647][14] = 1;
        layer_1_weights[648][14] = -1;
        layer_1_weights[649][14] = 1;
        layer_1_weights[650][14] = 1;
        layer_1_weights[651][14] = 1;
        layer_1_weights[652][14] = 2;
        layer_1_weights[653][14] = 1;
        layer_1_weights[654][14] = 1;
        layer_1_weights[655][14] = 2;
        layer_1_weights[656][14] = 1;
        layer_1_weights[657][14] = 0;
        layer_1_weights[658][14] = 1;
        layer_1_weights[659][14] = 1;
        layer_1_weights[660][14] = -1;
        layer_1_weights[661][14] = 1;
        layer_1_weights[662][14] = 2;
        layer_1_weights[663][14] = 1;
        layer_1_weights[664][14] = 2;
        layer_1_weights[665][14] = 3;
        layer_1_weights[666][14] = 4;
        layer_1_weights[667][14] = 1;
        layer_1_weights[668][14] = -1;
        layer_1_weights[669][14] = -1;
        layer_1_weights[670][14] = -3;
        layer_1_weights[671][14] = 1;
        layer_1_weights[672][14] = 0;
        layer_1_weights[673][14] = 0;
        layer_1_weights[674][14] = -2;
        layer_1_weights[675][14] = -6;
        layer_1_weights[676][14] = -4;
        layer_1_weights[677][14] = -5;
        layer_1_weights[678][14] = -2;
        layer_1_weights[679][14] = -2;
        layer_1_weights[680][14] = 0;
        layer_1_weights[681][14] = 0;
        layer_1_weights[682][14] = -1;
        layer_1_weights[683][14] = 0;
        layer_1_weights[684][14] = 1;
        layer_1_weights[685][14] = 1;
        layer_1_weights[686][14] = 0;
        layer_1_weights[687][14] = -1;
        layer_1_weights[688][14] = 0;
        layer_1_weights[689][14] = 0;
        layer_1_weights[690][14] = 2;
        layer_1_weights[691][14] = 2;
        layer_1_weights[692][14] = 2;
        layer_1_weights[693][14] = 1;
        layer_1_weights[694][14] = 0;
        layer_1_weights[695][14] = 1;
        layer_1_weights[696][14] = -1;
        layer_1_weights[697][14] = 4;
        layer_1_weights[698][14] = 2;
        layer_1_weights[699][14] = 1;
        layer_1_weights[700][14] = 0;
        layer_1_weights[701][14] = 0;
        layer_1_weights[702][14] = 0;
        layer_1_weights[703][14] = -5;
        layer_1_weights[704][14] = -3;
        layer_1_weights[705][14] = -3;
        layer_1_weights[706][14] = -2;
        layer_1_weights[707][14] = -2;
        layer_1_weights[708][14] = -3;
        layer_1_weights[709][14] = -3;
        layer_1_weights[710][14] = -3;
        layer_1_weights[711][14] = -2;
        layer_1_weights[712][14] = -2;
        layer_1_weights[713][14] = -1;
        layer_1_weights[714][14] = 0;
        layer_1_weights[715][14] = 0;
        layer_1_weights[716][14] = -2;
        layer_1_weights[717][14] = -1;
        layer_1_weights[718][14] = 0;
        layer_1_weights[719][14] = -1;
        layer_1_weights[720][14] = -1;
        layer_1_weights[721][14] = -2;
        layer_1_weights[722][14] = -3;
        layer_1_weights[723][14] = -2;
        layer_1_weights[724][14] = -5;
        layer_1_weights[725][14] = 3;
        layer_1_weights[726][14] = 1;
        layer_1_weights[727][14] = -1;
        layer_1_weights[728][14] = 0;
        layer_1_weights[729][14] = 0;
        layer_1_weights[730][14] = 0;
        layer_1_weights[731][14] = 2;
        layer_1_weights[732][14] = 2;
        layer_1_weights[733][14] = 1;
        layer_1_weights[734][14] = 1;
        layer_1_weights[735][14] = 0;
        layer_1_weights[736][14] = -1;
        layer_1_weights[737][14] = -1;
        layer_1_weights[738][14] = -3;
        layer_1_weights[739][14] = -1;
        layer_1_weights[740][14] = 1;
        layer_1_weights[741][14] = 0;
        layer_1_weights[742][14] = -1;
        layer_1_weights[743][14] = -3;
        layer_1_weights[744][14] = -5;
        layer_1_weights[745][14] = -4;
        layer_1_weights[746][14] = -5;
        layer_1_weights[747][14] = -3;
        layer_1_weights[748][14] = -4;
        layer_1_weights[749][14] = -2;
        layer_1_weights[750][14] = -2;
        layer_1_weights[751][14] = 1;
        layer_1_weights[752][14] = -1;
        layer_1_weights[753][14] = -2;
        layer_1_weights[754][14] = 1;
        layer_1_weights[755][14] = 0;
        layer_1_weights[756][14] = -1;
        layer_1_weights[757][14] = 0;
        layer_1_weights[758][14] = 0;
        layer_1_weights[759][14] = 0;
        layer_1_weights[760][14] = -3;
        layer_1_weights[761][14] = -4;
        layer_1_weights[762][14] = 2;
        layer_1_weights[763][14] = 2;
        layer_1_weights[764][14] = 1;
        layer_1_weights[765][14] = 3;
        layer_1_weights[766][14] = 1;
        layer_1_weights[767][14] = 1;
        layer_1_weights[768][14] = 1;
        layer_1_weights[769][14] = 0;
        layer_1_weights[770][14] = -1;
        layer_1_weights[771][14] = -1;
        layer_1_weights[772][14] = -2;
        layer_1_weights[773][14] = 0;
        layer_1_weights[774][14] = 1;
        layer_1_weights[775][14] = 0;
        layer_1_weights[776][14] = 1;
        layer_1_weights[777][14] = -2;
        layer_1_weights[778][14] = -2;
        layer_1_weights[779][14] = -3;
        layer_1_weights[780][14] = 0;
        layer_1_weights[781][14] = 1;
        layer_1_weights[782][14] = 0;
        layer_1_weights[783][14] = -1;
        layer_1_weights[0][15] = 0;
        layer_1_weights[1][15] = 0;
        layer_1_weights[2][15] = 0;
        layer_1_weights[3][15] = 0;
        layer_1_weights[4][15] = 0;
        layer_1_weights[5][15] = 1;
        layer_1_weights[6][15] = 0;
        layer_1_weights[7][15] = 0;
        layer_1_weights[8][15] = 1;
        layer_1_weights[9][15] = 0;
        layer_1_weights[10][15] = 0;
        layer_1_weights[11][15] = 1;
        layer_1_weights[12][15] = 0;
        layer_1_weights[13][15] = -1;
        layer_1_weights[14][15] = 0;
        layer_1_weights[15][15] = 0;
        layer_1_weights[16][15] = 0;
        layer_1_weights[17][15] = 0;
        layer_1_weights[18][15] = 0;
        layer_1_weights[19][15] = 1;
        layer_1_weights[20][15] = 0;
        layer_1_weights[21][15] = 0;
        layer_1_weights[22][15] = 0;
        layer_1_weights[23][15] = 0;
        layer_1_weights[24][15] = 0;
        layer_1_weights[25][15] = 0;
        layer_1_weights[26][15] = 0;
        layer_1_weights[27][15] = -1;
        layer_1_weights[28][15] = 0;
        layer_1_weights[29][15] = 0;
        layer_1_weights[30][15] = -1;
        layer_1_weights[31][15] = 0;
        layer_1_weights[32][15] = -1;
        layer_1_weights[33][15] = 0;
        layer_1_weights[34][15] = 0;
        layer_1_weights[35][15] = 0;
        layer_1_weights[36][15] = -1;
        layer_1_weights[37][15] = 1;
        layer_1_weights[38][15] = 0;
        layer_1_weights[39][15] = 3;
        layer_1_weights[40][15] = 2;
        layer_1_weights[41][15] = 1;
        layer_1_weights[42][15] = 0;
        layer_1_weights[43][15] = -1;
        layer_1_weights[44][15] = -2;
        layer_1_weights[45][15] = 0;
        layer_1_weights[46][15] = 2;
        layer_1_weights[47][15] = 1;
        layer_1_weights[48][15] = -3;
        layer_1_weights[49][15] = 0;
        layer_1_weights[50][15] = -2;
        layer_1_weights[51][15] = -1;
        layer_1_weights[52][15] = 0;
        layer_1_weights[53][15] = 0;
        layer_1_weights[54][15] = -1;
        layer_1_weights[55][15] = 1;
        layer_1_weights[56][15] = 0;
        layer_1_weights[57][15] = 0;
        layer_1_weights[58][15] = 0;
        layer_1_weights[59][15] = 0;
        layer_1_weights[60][15] = -2;
        layer_1_weights[61][15] = 1;
        layer_1_weights[62][15] = 0;
        layer_1_weights[63][15] = 0;
        layer_1_weights[64][15] = -1;
        layer_1_weights[65][15] = -3;
        layer_1_weights[66][15] = -3;
        layer_1_weights[67][15] = -4;
        layer_1_weights[68][15] = -1;
        layer_1_weights[69][15] = -5;
        layer_1_weights[70][15] = -7;
        layer_1_weights[71][15] = -2;
        layer_1_weights[72][15] = -4;
        layer_1_weights[73][15] = -5;
        layer_1_weights[74][15] = -6;
        layer_1_weights[75][15] = 4;
        layer_1_weights[76][15] = 0;
        layer_1_weights[77][15] = 3;
        layer_1_weights[78][15] = 2;
        layer_1_weights[79][15] = 2;
        layer_1_weights[80][15] = 2;
        layer_1_weights[81][15] = -1;
        layer_1_weights[82][15] = 0;
        layer_1_weights[83][15] = 0;
        layer_1_weights[84][15] = 0;
        layer_1_weights[85][15] = -1;
        layer_1_weights[86][15] = 2;
        layer_1_weights[87][15] = 1;
        layer_1_weights[88][15] = 0;
        layer_1_weights[89][15] = -2;
        layer_1_weights[90][15] = -2;
        layer_1_weights[91][15] = -1;
        layer_1_weights[92][15] = -4;
        layer_1_weights[93][15] = -5;
        layer_1_weights[94][15] = -5;
        layer_1_weights[95][15] = -6;
        layer_1_weights[96][15] = -4;
        layer_1_weights[97][15] = -7;
        layer_1_weights[98][15] = -6;
        layer_1_weights[99][15] = -8;
        layer_1_weights[100][15] = -5;
        layer_1_weights[101][15] = -3;
        layer_1_weights[102][15] = 0;
        layer_1_weights[103][15] = 0;
        layer_1_weights[104][15] = 0;
        layer_1_weights[105][15] = -3;
        layer_1_weights[106][15] = -1;
        layer_1_weights[107][15] = 1;
        layer_1_weights[108][15] = -2;
        layer_1_weights[109][15] = 0;
        layer_1_weights[110][15] = 1;
        layer_1_weights[111][15] = 0;
        layer_1_weights[112][15] = 0;
        layer_1_weights[113][15] = 1;
        layer_1_weights[114][15] = 3;
        layer_1_weights[115][15] = 3;
        layer_1_weights[116][15] = 2;
        layer_1_weights[117][15] = -2;
        layer_1_weights[118][15] = -2;
        layer_1_weights[119][15] = -2;
        layer_1_weights[120][15] = -2;
        layer_1_weights[121][15] = -2;
        layer_1_weights[122][15] = -3;
        layer_1_weights[123][15] = -3;
        layer_1_weights[124][15] = -1;
        layer_1_weights[125][15] = -2;
        layer_1_weights[126][15] = -2;
        layer_1_weights[127][15] = -2;
        layer_1_weights[128][15] = -1;
        layer_1_weights[129][15] = -2;
        layer_1_weights[130][15] = 0;
        layer_1_weights[131][15] = 2;
        layer_1_weights[132][15] = 1;
        layer_1_weights[133][15] = 1;
        layer_1_weights[134][15] = 0;
        layer_1_weights[135][15] = 0;
        layer_1_weights[136][15] = -1;
        layer_1_weights[137][15] = -6;
        layer_1_weights[138][15] = -1;
        layer_1_weights[139][15] = 1;
        layer_1_weights[140][15] = 0;
        layer_1_weights[141][15] = 0;
        layer_1_weights[142][15] = 0;
        layer_1_weights[143][15] = 3;
        layer_1_weights[144][15] = -1;
        layer_1_weights[145][15] = 1;
        layer_1_weights[146][15] = -1;
        layer_1_weights[147][15] = 2;
        layer_1_weights[148][15] = -1;
        layer_1_weights[149][15] = -3;
        layer_1_weights[150][15] = -1;
        layer_1_weights[151][15] = -1;
        layer_1_weights[152][15] = -1;
        layer_1_weights[153][15] = 0;
        layer_1_weights[154][15] = 0;
        layer_1_weights[155][15] = 0;
        layer_1_weights[156][15] = -1;
        layer_1_weights[157][15] = 0;
        layer_1_weights[158][15] = -2;
        layer_1_weights[159][15] = -1;
        layer_1_weights[160][15] = -2;
        layer_1_weights[161][15] = 0;
        layer_1_weights[162][15] = 1;
        layer_1_weights[163][15] = -1;
        layer_1_weights[164][15] = 2;
        layer_1_weights[165][15] = -3;
        layer_1_weights[166][15] = 0;
        layer_1_weights[167][15] = 2;
        layer_1_weights[168][15] = 0;
        layer_1_weights[169][15] = 0;
        layer_1_weights[170][15] = -1;
        layer_1_weights[171][15] = 2;
        layer_1_weights[172][15] = -1;
        layer_1_weights[173][15] = 0;
        layer_1_weights[174][15] = -2;
        layer_1_weights[175][15] = 2;
        layer_1_weights[176][15] = 0;
        layer_1_weights[177][15] = 0;
        layer_1_weights[178][15] = 0;
        layer_1_weights[179][15] = 0;
        layer_1_weights[180][15] = -1;
        layer_1_weights[181][15] = 0;
        layer_1_weights[182][15] = 0;
        layer_1_weights[183][15] = 0;
        layer_1_weights[184][15] = 0;
        layer_1_weights[185][15] = 0;
        layer_1_weights[186][15] = -1;
        layer_1_weights[187][15] = 0;
        layer_1_weights[188][15] = -2;
        layer_1_weights[189][15] = 1;
        layer_1_weights[190][15] = 0;
        layer_1_weights[191][15] = 1;
        layer_1_weights[192][15] = 0;
        layer_1_weights[193][15] = -3;
        layer_1_weights[194][15] = -1;
        layer_1_weights[195][15] = 2;
        layer_1_weights[196][15] = 1;
        layer_1_weights[197][15] = -4;
        layer_1_weights[198][15] = 0;
        layer_1_weights[199][15] = 0;
        layer_1_weights[200][15] = 2;
        layer_1_weights[201][15] = -1;
        layer_1_weights[202][15] = 1;
        layer_1_weights[203][15] = -1;
        layer_1_weights[204][15] = 0;
        layer_1_weights[205][15] = 1;
        layer_1_weights[206][15] = 0;
        layer_1_weights[207][15] = -1;
        layer_1_weights[208][15] = 2;
        layer_1_weights[209][15] = 0;
        layer_1_weights[210][15] = -1;
        layer_1_weights[211][15] = -1;
        layer_1_weights[212][15] = -1;
        layer_1_weights[213][15] = 2;
        layer_1_weights[214][15] = 1;
        layer_1_weights[215][15] = 0;
        layer_1_weights[216][15] = 1;
        layer_1_weights[217][15] = 0;
        layer_1_weights[218][15] = -1;
        layer_1_weights[219][15] = 1;
        layer_1_weights[220][15] = -3;
        layer_1_weights[221][15] = -2;
        layer_1_weights[222][15] = 1;
        layer_1_weights[223][15] = 2;
        layer_1_weights[224][15] = 2;
        layer_1_weights[225][15] = -2;
        layer_1_weights[226][15] = 3;
        layer_1_weights[227][15] = 1;
        layer_1_weights[228][15] = 3;
        layer_1_weights[229][15] = -3;
        layer_1_weights[230][15] = 0;
        layer_1_weights[231][15] = -1;
        layer_1_weights[232][15] = 0;
        layer_1_weights[233][15] = -1;
        layer_1_weights[234][15] = 1;
        layer_1_weights[235][15] = 0;
        layer_1_weights[236][15] = 0;
        layer_1_weights[237][15] = 0;
        layer_1_weights[238][15] = 2;
        layer_1_weights[239][15] = 2;
        layer_1_weights[240][15] = 1;
        layer_1_weights[241][15] = 0;
        layer_1_weights[242][15] = -1;
        layer_1_weights[243][15] = 0;
        layer_1_weights[244][15] = 0;
        layer_1_weights[245][15] = 0;
        layer_1_weights[246][15] = -1;
        layer_1_weights[247][15] = -3;
        layer_1_weights[248][15] = -6;
        layer_1_weights[249][15] = -3;
        layer_1_weights[250][15] = 0;
        layer_1_weights[251][15] = -4;
        layer_1_weights[252][15] = 0;
        layer_1_weights[253][15] = 2;
        layer_1_weights[254][15] = 2;
        layer_1_weights[255][15] = -4;
        layer_1_weights[256][15] = -2;
        layer_1_weights[257][15] = -1;
        layer_1_weights[258][15] = 1;
        layer_1_weights[259][15] = 0;
        layer_1_weights[260][15] = 1;
        layer_1_weights[261][15] = 0;
        layer_1_weights[262][15] = 0;
        layer_1_weights[263][15] = 0;
        layer_1_weights[264][15] = -1;
        layer_1_weights[265][15] = 1;
        layer_1_weights[266][15] = 2;
        layer_1_weights[267][15] = 1;
        layer_1_weights[268][15] = 1;
        layer_1_weights[269][15] = 0;
        layer_1_weights[270][15] = 0;
        layer_1_weights[271][15] = 1;
        layer_1_weights[272][15] = -1;
        layer_1_weights[273][15] = 0;
        layer_1_weights[274][15] = 0;
        layer_1_weights[275][15] = -3;
        layer_1_weights[276][15] = -4;
        layer_1_weights[277][15] = -1;
        layer_1_weights[278][15] = -1;
        layer_1_weights[279][15] = 2;
        layer_1_weights[280][15] = 1;
        layer_1_weights[281][15] = 5;
        layer_1_weights[282][15] = 2;
        layer_1_weights[283][15] = -2;
        layer_1_weights[284][15] = 1;
        layer_1_weights[285][15] = -1;
        layer_1_weights[286][15] = -2;
        layer_1_weights[287][15] = -1;
        layer_1_weights[288][15] = -1;
        layer_1_weights[289][15] = 0;
        layer_1_weights[290][15] = -2;
        layer_1_weights[291][15] = -2;
        layer_1_weights[292][15] = -1;
        layer_1_weights[293][15] = 1;
        layer_1_weights[294][15] = 3;
        layer_1_weights[295][15] = 1;
        layer_1_weights[296][15] = 2;
        layer_1_weights[297][15] = 1;
        layer_1_weights[298][15] = 0;
        layer_1_weights[299][15] = 1;
        layer_1_weights[300][15] = -1;
        layer_1_weights[301][15] = -2;
        layer_1_weights[302][15] = -1;
        layer_1_weights[303][15] = -2;
        layer_1_weights[304][15] = -6;
        layer_1_weights[305][15] = -3;
        layer_1_weights[306][15] = 0;
        layer_1_weights[307][15] = 3;
        layer_1_weights[308][15] = 3;
        layer_1_weights[309][15] = 5;
        layer_1_weights[310][15] = 0;
        layer_1_weights[311][15] = 1;
        layer_1_weights[312][15] = -2;
        layer_1_weights[313][15] = 0;
        layer_1_weights[314][15] = -2;
        layer_1_weights[315][15] = -1;
        layer_1_weights[316][15] = -1;
        layer_1_weights[317][15] = -1;
        layer_1_weights[318][15] = 0;
        layer_1_weights[319][15] = 1;
        layer_1_weights[320][15] = 0;
        layer_1_weights[321][15] = 1;
        layer_1_weights[322][15] = 2;
        layer_1_weights[323][15] = 2;
        layer_1_weights[324][15] = 1;
        layer_1_weights[325][15] = 1;
        layer_1_weights[326][15] = 2;
        layer_1_weights[327][15] = 0;
        layer_1_weights[328][15] = 0;
        layer_1_weights[329][15] = -1;
        layer_1_weights[330][15] = -1;
        layer_1_weights[331][15] = -4;
        layer_1_weights[332][15] = -4;
        layer_1_weights[333][15] = -6;
        layer_1_weights[334][15] = -1;
        layer_1_weights[335][15] = -2;
        layer_1_weights[336][15] = 1;
        layer_1_weights[337][15] = 5;
        layer_1_weights[338][15] = 3;
        layer_1_weights[339][15] = 1;
        layer_1_weights[340][15] = -3;
        layer_1_weights[341][15] = -3;
        layer_1_weights[342][15] = 0;
        layer_1_weights[343][15] = 1;
        layer_1_weights[344][15] = 0;
        layer_1_weights[345][15] = 0;
        layer_1_weights[346][15] = 0;
        layer_1_weights[347][15] = 1;
        layer_1_weights[348][15] = 1;
        layer_1_weights[349][15] = 2;
        layer_1_weights[350][15] = 1;
        layer_1_weights[351][15] = 3;
        layer_1_weights[352][15] = 2;
        layer_1_weights[353][15] = 2;
        layer_1_weights[354][15] = 2;
        layer_1_weights[355][15] = 0;
        layer_1_weights[356][15] = 1;
        layer_1_weights[357][15] = 0;
        layer_1_weights[358][15] = -2;
        layer_1_weights[359][15] = -6;
        layer_1_weights[360][15] = -4;
        layer_1_weights[361][15] = -4;
        layer_1_weights[362][15] = -3;
        layer_1_weights[363][15] = 3;
        layer_1_weights[364][15] = -1;
        layer_1_weights[365][15] = 2;
        layer_1_weights[366][15] = 5;
        layer_1_weights[367][15] = 1;
        layer_1_weights[368][15] = -1;
        layer_1_weights[369][15] = -3;
        layer_1_weights[370][15] = 0;
        layer_1_weights[371][15] = 0;
        layer_1_weights[372][15] = 0;
        layer_1_weights[373][15] = 0;
        layer_1_weights[374][15] = 0;
        layer_1_weights[375][15] = 2;
        layer_1_weights[376][15] = 2;
        layer_1_weights[377][15] = 1;
        layer_1_weights[378][15] = 2;
        layer_1_weights[379][15] = 1;
        layer_1_weights[380][15] = 0;
        layer_1_weights[381][15] = 2;
        layer_1_weights[382][15] = 1;
        layer_1_weights[383][15] = 2;
        layer_1_weights[384][15] = 2;
        layer_1_weights[385][15] = 1;
        layer_1_weights[386][15] = -3;
        layer_1_weights[387][15] = -4;
        layer_1_weights[388][15] = -7;
        layer_1_weights[389][15] = -4;
        layer_1_weights[390][15] = -6;
        layer_1_weights[391][15] = 0;
        layer_1_weights[392][15] = -2;
        layer_1_weights[393][15] = 1;
        layer_1_weights[394][15] = 4;
        layer_1_weights[395][15] = 2;
        layer_1_weights[396][15] = 2;
        layer_1_weights[397][15] = 0;
        layer_1_weights[398][15] = -3;
        layer_1_weights[399][15] = -2;
        layer_1_weights[400][15] = -1;
        layer_1_weights[401][15] = 0;
        layer_1_weights[402][15] = 0;
        layer_1_weights[403][15] = 3;
        layer_1_weights[404][15] = 2;
        layer_1_weights[405][15] = 2;
        layer_1_weights[406][15] = 1;
        layer_1_weights[407][15] = 1;
        layer_1_weights[408][15] = 2;
        layer_1_weights[409][15] = 2;
        layer_1_weights[410][15] = 2;
        layer_1_weights[411][15] = 2;
        layer_1_weights[412][15] = 2;
        layer_1_weights[413][15] = -1;
        layer_1_weights[414][15] = -1;
        layer_1_weights[415][15] = -4;
        layer_1_weights[416][15] = -5;
        layer_1_weights[417][15] = -4;
        layer_1_weights[418][15] = -5;
        layer_1_weights[419][15] = 0;
        layer_1_weights[420][15] = -2;
        layer_1_weights[421][15] = 0;
        layer_1_weights[422][15] = 0;
        layer_1_weights[423][15] = 2;
        layer_1_weights[424][15] = -2;
        layer_1_weights[425][15] = -3;
        layer_1_weights[426][15] = -1;
        layer_1_weights[427][15] = -3;
        layer_1_weights[428][15] = -3;
        layer_1_weights[429][15] = 0;
        layer_1_weights[430][15] = 1;
        layer_1_weights[431][15] = 1;
        layer_1_weights[432][15] = 2;
        layer_1_weights[433][15] = 2;
        layer_1_weights[434][15] = 0;
        layer_1_weights[435][15] = 2;
        layer_1_weights[436][15] = 1;
        layer_1_weights[437][15] = 1;
        layer_1_weights[438][15] = 3;
        layer_1_weights[439][15] = 1;
        layer_1_weights[440][15] = 0;
        layer_1_weights[441][15] = -4;
        layer_1_weights[442][15] = -3;
        layer_1_weights[443][15] = -3;
        layer_1_weights[444][15] = -3;
        layer_1_weights[445][15] = -5;
        layer_1_weights[446][15] = -3;
        layer_1_weights[447][15] = 0;
        layer_1_weights[448][15] = 2;
        layer_1_weights[449][15] = -3;
        layer_1_weights[450][15] = -2;
        layer_1_weights[451][15] = -2;
        layer_1_weights[452][15] = 2;
        layer_1_weights[453][15] = -2;
        layer_1_weights[454][15] = -3;
        layer_1_weights[455][15] = -3;
        layer_1_weights[456][15] = -2;
        layer_1_weights[457][15] = 0;
        layer_1_weights[458][15] = 0;
        layer_1_weights[459][15] = 2;
        layer_1_weights[460][15] = 2;
        layer_1_weights[461][15] = 2;
        layer_1_weights[462][15] = 1;
        layer_1_weights[463][15] = 0;
        layer_1_weights[464][15] = 1;
        layer_1_weights[465][15] = 3;
        layer_1_weights[466][15] = 1;
        layer_1_weights[467][15] = 1;
        layer_1_weights[468][15] = -1;
        layer_1_weights[469][15] = -3;
        layer_1_weights[470][15] = -5;
        layer_1_weights[471][15] = -6;
        layer_1_weights[472][15] = -4;
        layer_1_weights[473][15] = -5;
        layer_1_weights[474][15] = -3;
        layer_1_weights[475][15] = -3;
        layer_1_weights[476][15] = 0;
        layer_1_weights[477][15] = 1;
        layer_1_weights[478][15] = -2;
        layer_1_weights[479][15] = -1;
        layer_1_weights[480][15] = 1;
        layer_1_weights[481][15] = -2;
        layer_1_weights[482][15] = -1;
        layer_1_weights[483][15] = -4;
        layer_1_weights[484][15] = -1;
        layer_1_weights[485][15] = -1;
        layer_1_weights[486][15] = 0;
        layer_1_weights[487][15] = 0;
        layer_1_weights[488][15] = 1;
        layer_1_weights[489][15] = 1;
        layer_1_weights[490][15] = 0;
        layer_1_weights[491][15] = 0;
        layer_1_weights[492][15] = 2;
        layer_1_weights[493][15] = 0;
        layer_1_weights[494][15] = 1;
        layer_1_weights[495][15] = 0;
        layer_1_weights[496][15] = -3;
        layer_1_weights[497][15] = -4;
        layer_1_weights[498][15] = -3;
        layer_1_weights[499][15] = -3;
        layer_1_weights[500][15] = -2;
        layer_1_weights[501][15] = 1;
        layer_1_weights[502][15] = 0;
        layer_1_weights[503][15] = -3;
        layer_1_weights[504][15] = -2;
        layer_1_weights[505][15] = 1;
        layer_1_weights[506][15] = -3;
        layer_1_weights[507][15] = 0;
        layer_1_weights[508][15] = -2;
        layer_1_weights[509][15] = -3;
        layer_1_weights[510][15] = -2;
        layer_1_weights[511][15] = -1;
        layer_1_weights[512][15] = -3;
        layer_1_weights[513][15] = 0;
        layer_1_weights[514][15] = 0;
        layer_1_weights[515][15] = 1;
        layer_1_weights[516][15] = 1;
        layer_1_weights[517][15] = 0;
        layer_1_weights[518][15] = 1;
        layer_1_weights[519][15] = 0;
        layer_1_weights[520][15] = -1;
        layer_1_weights[521][15] = -1;
        layer_1_weights[522][15] = 0;
        layer_1_weights[523][15] = -2;
        layer_1_weights[524][15] = -3;
        layer_1_weights[525][15] = -2;
        layer_1_weights[526][15] = -4;
        layer_1_weights[527][15] = -4;
        layer_1_weights[528][15] = -5;
        layer_1_weights[529][15] = 1;
        layer_1_weights[530][15] = 3;
        layer_1_weights[531][15] = 3;
        layer_1_weights[532][15] = 0;
        layer_1_weights[533][15] = -1;
        layer_1_weights[534][15] = -1;
        layer_1_weights[535][15] = 1;
        layer_1_weights[536][15] = -1;
        layer_1_weights[537][15] = -2;
        layer_1_weights[538][15] = -2;
        layer_1_weights[539][15] = 0;
        layer_1_weights[540][15] = -2;
        layer_1_weights[541][15] = -2;
        layer_1_weights[542][15] = 0;
        layer_1_weights[543][15] = 1;
        layer_1_weights[544][15] = 1;
        layer_1_weights[545][15] = 0;
        layer_1_weights[546][15] = 0;
        layer_1_weights[547][15] = 0;
        layer_1_weights[548][15] = -1;
        layer_1_weights[549][15] = -1;
        layer_1_weights[550][15] = 0;
        layer_1_weights[551][15] = -2;
        layer_1_weights[552][15] = -3;
        layer_1_weights[553][15] = -2;
        layer_1_weights[554][15] = -4;
        layer_1_weights[555][15] = -3;
        layer_1_weights[556][15] = -3;
        layer_1_weights[557][15] = 1;
        layer_1_weights[558][15] = 1;
        layer_1_weights[559][15] = 2;
        layer_1_weights[560][15] = 0;
        layer_1_weights[561][15] = 3;
        layer_1_weights[562][15] = -2;
        layer_1_weights[563][15] = -2;
        layer_1_weights[564][15] = 0;
        layer_1_weights[565][15] = 0;
        layer_1_weights[566][15] = 0;
        layer_1_weights[567][15] = -2;
        layer_1_weights[568][15] = -2;
        layer_1_weights[569][15] = -1;
        layer_1_weights[570][15] = 0;
        layer_1_weights[571][15] = 0;
        layer_1_weights[572][15] = 0;
        layer_1_weights[573][15] = 0;
        layer_1_weights[574][15] = 0;
        layer_1_weights[575][15] = -1;
        layer_1_weights[576][15] = -1;
        layer_1_weights[577][15] = -2;
        layer_1_weights[578][15] = -2;
        layer_1_weights[579][15] = -2;
        layer_1_weights[580][15] = -2;
        layer_1_weights[581][15] = 0;
        layer_1_weights[582][15] = -1;
        layer_1_weights[583][15] = -3;
        layer_1_weights[584][15] = -1;
        layer_1_weights[585][15] = -1;
        layer_1_weights[586][15] = 1;
        layer_1_weights[587][15] = 2;
        layer_1_weights[588][15] = 0;
        layer_1_weights[589][15] = -3;
        layer_1_weights[590][15] = -2;
        layer_1_weights[591][15] = -3;
        layer_1_weights[592][15] = -3;
        layer_1_weights[593][15] = -1;
        layer_1_weights[594][15] = 0;
        layer_1_weights[595][15] = -1;
        layer_1_weights[596][15] = -1;
        layer_1_weights[597][15] = -1;
        layer_1_weights[598][15] = 1;
        layer_1_weights[599][15] = 1;
        layer_1_weights[600][15] = 0;
        layer_1_weights[601][15] = -2;
        layer_1_weights[602][15] = -1;
        layer_1_weights[603][15] = -1;
        layer_1_weights[604][15] = -1;
        layer_1_weights[605][15] = -1;
        layer_1_weights[606][15] = -1;
        layer_1_weights[607][15] = -1;
        layer_1_weights[608][15] = -2;
        layer_1_weights[609][15] = -5;
        layer_1_weights[610][15] = -1;
        layer_1_weights[611][15] = -1;
        layer_1_weights[612][15] = 0;
        layer_1_weights[613][15] = -2;
        layer_1_weights[614][15] = 0;
        layer_1_weights[615][15] = 0;
        layer_1_weights[616][15] = 0;
        layer_1_weights[617][15] = 1;
        layer_1_weights[618][15] = -3;
        layer_1_weights[619][15] = -1;
        layer_1_weights[620][15] = -2;
        layer_1_weights[621][15] = 0;
        layer_1_weights[622][15] = 1;
        layer_1_weights[623][15] = 1;
        layer_1_weights[624][15] = 1;
        layer_1_weights[625][15] = 0;
        layer_1_weights[626][15] = 1;
        layer_1_weights[627][15] = -1;
        layer_1_weights[628][15] = -1;
        layer_1_weights[629][15] = -1;
        layer_1_weights[630][15] = 0;
        layer_1_weights[631][15] = 1;
        layer_1_weights[632][15] = -1;
        layer_1_weights[633][15] = -1;
        layer_1_weights[634][15] = -1;
        layer_1_weights[635][15] = -1;
        layer_1_weights[636][15] = -3;
        layer_1_weights[637][15] = -2;
        layer_1_weights[638][15] = -3;
        layer_1_weights[639][15] = 1;
        layer_1_weights[640][15] = 2;
        layer_1_weights[641][15] = -1;
        layer_1_weights[642][15] = 3;
        layer_1_weights[643][15] = 0;
        layer_1_weights[644][15] = 0;
        layer_1_weights[645][15] = 0;
        layer_1_weights[646][15] = -4;
        layer_1_weights[647][15] = -3;
        layer_1_weights[648][15] = -4;
        layer_1_weights[649][15] = 0;
        layer_1_weights[650][15] = 0;
        layer_1_weights[651][15] = 1;
        layer_1_weights[652][15] = 0;
        layer_1_weights[653][15] = 1;
        layer_1_weights[654][15] = 1;
        layer_1_weights[655][15] = -1;
        layer_1_weights[656][15] = 1;
        layer_1_weights[657][15] = 0;
        layer_1_weights[658][15] = 0;
        layer_1_weights[659][15] = 0;
        layer_1_weights[660][15] = -1;
        layer_1_weights[661][15] = 0;
        layer_1_weights[662][15] = -1;
        layer_1_weights[663][15] = -3;
        layer_1_weights[664][15] = -3;
        layer_1_weights[665][15] = -5;
        layer_1_weights[666][15] = 1;
        layer_1_weights[667][15] = 0;
        layer_1_weights[668][15] = 0;
        layer_1_weights[669][15] = -1;
        layer_1_weights[670][15] = 3;
        layer_1_weights[671][15] = -1;
        layer_1_weights[672][15] = 1;
        layer_1_weights[673][15] = -1;
        layer_1_weights[674][15] = -2;
        layer_1_weights[675][15] = -3;
        layer_1_weights[676][15] = -1;
        layer_1_weights[677][15] = 2;
        layer_1_weights[678][15] = 0;
        layer_1_weights[679][15] = 2;
        layer_1_weights[680][15] = -2;
        layer_1_weights[681][15] = 0;
        layer_1_weights[682][15] = -2;
        layer_1_weights[683][15] = -2;
        layer_1_weights[684][15] = -1;
        layer_1_weights[685][15] = -1;
        layer_1_weights[686][15] = -2;
        layer_1_weights[687][15] = -1;
        layer_1_weights[688][15] = -2;
        layer_1_weights[689][15] = -2;
        layer_1_weights[690][15] = 2;
        layer_1_weights[691][15] = -3;
        layer_1_weights[692][15] = 0;
        layer_1_weights[693][15] = -1;
        layer_1_weights[694][15] = 0;
        layer_1_weights[695][15] = 2;
        layer_1_weights[696][15] = -3;
        layer_1_weights[697][15] = 1;
        layer_1_weights[698][15] = -1;
        layer_1_weights[699][15] = -1;
        layer_1_weights[700][15] = 0;
        layer_1_weights[701][15] = 0;
        layer_1_weights[702][15] = 0;
        layer_1_weights[703][15] = 3;
        layer_1_weights[704][15] = 3;
        layer_1_weights[705][15] = 0;
        layer_1_weights[706][15] = 0;
        layer_1_weights[707][15] = 0;
        layer_1_weights[708][15] = -1;
        layer_1_weights[709][15] = 0;
        layer_1_weights[710][15] = -1;
        layer_1_weights[711][15] = -2;
        layer_1_weights[712][15] = -1;
        layer_1_weights[713][15] = -2;
        layer_1_weights[714][15] = -1;
        layer_1_weights[715][15] = -2;
        layer_1_weights[716][15] = -3;
        layer_1_weights[717][15] = -3;
        layer_1_weights[718][15] = -1;
        layer_1_weights[719][15] = 1;
        layer_1_weights[720][15] = -2;
        layer_1_weights[721][15] = -1;
        layer_1_weights[722][15] = -1;
        layer_1_weights[723][15] = 5;
        layer_1_weights[724][15] = 3;
        layer_1_weights[725][15] = -3;
        layer_1_weights[726][15] = -2;
        layer_1_weights[727][15] = 0;
        layer_1_weights[728][15] = 0;
        layer_1_weights[729][15] = 0;
        layer_1_weights[730][15] = 0;
        layer_1_weights[731][15] = -2;
        layer_1_weights[732][15] = 1;
        layer_1_weights[733][15] = 1;
        layer_1_weights[734][15] = 1;
        layer_1_weights[735][15] = 4;
        layer_1_weights[736][15] = 0;
        layer_1_weights[737][15] = 0;
        layer_1_weights[738][15] = -2;
        layer_1_weights[739][15] = -1;
        layer_1_weights[740][15] = 0;
        layer_1_weights[741][15] = 0;
        layer_1_weights[742][15] = 1;
        layer_1_weights[743][15] = -1;
        layer_1_weights[744][15] = 0;
        layer_1_weights[745][15] = -1;
        layer_1_weights[746][15] = -1;
        layer_1_weights[747][15] = -1;
        layer_1_weights[748][15] = -2;
        layer_1_weights[749][15] = -2;
        layer_1_weights[750][15] = -3;
        layer_1_weights[751][15] = -2;
        layer_1_weights[752][15] = 0;
        layer_1_weights[753][15] = 2;
        layer_1_weights[754][15] = 0;
        layer_1_weights[755][15] = 0;
        layer_1_weights[756][15] = 0;
        layer_1_weights[757][15] = 0;
        layer_1_weights[758][15] = 1;
        layer_1_weights[759][15] = 0;
        layer_1_weights[760][15] = 2;
        layer_1_weights[761][15] = 3;
        layer_1_weights[762][15] = -2;
        layer_1_weights[763][15] = -2;
        layer_1_weights[764][15] = -1;
        layer_1_weights[765][15] = -2;
        layer_1_weights[766][15] = 1;
        layer_1_weights[767][15] = 1;
        layer_1_weights[768][15] = 1;
        layer_1_weights[769][15] = 3;
        layer_1_weights[770][15] = -4;
        layer_1_weights[771][15] = -3;
        layer_1_weights[772][15] = 0;
        layer_1_weights[773][15] = 1;
        layer_1_weights[774][15] = -2;
        layer_1_weights[775][15] = 0;
        layer_1_weights[776][15] = 2;
        layer_1_weights[777][15] = 0;
        layer_1_weights[778][15] = 0;
        layer_1_weights[779][15] = 0;
        layer_1_weights[780][15] = -1;
        layer_1_weights[781][15] = 0;
        layer_1_weights[782][15] = 0;
        layer_1_weights[783][15] = 1;
        layer_1_biases[0] = -1;
        layer_1_biases[1] = -1;
        layer_1_biases[2] = 3;
        layer_1_biases[3] = 6;
        layer_1_biases[4] = -2;
        layer_1_biases[5] = -3;
        layer_1_biases[6] = 6;
        layer_1_biases[7] = -2;
        layer_1_biases[8] = 0;
        layer_1_biases[9] = 7;
        layer_1_biases[10] = -2;
        layer_1_biases[11] = 1;
        layer_1_biases[12] = -1;
        layer_1_biases[13] = -4;
        layer_1_biases[14] = -5;
        layer_1_biases[15] = 1;
        layer_2_weights[0][0] = 0;
        layer_2_weights[1][0] = 0;
        layer_2_weights[2][0] = 2;
        layer_2_weights[3][0] = 0;
        layer_2_weights[4][0] = 2;
        layer_2_weights[5][0] = -6;
        layer_2_weights[6][0] = -2;
        layer_2_weights[7][0] = 1;
        layer_2_weights[8][0] = 3;
        layer_2_weights[9][0] = -9;
        layer_2_weights[10][0] = 5;
        layer_2_weights[11][0] = 0;
        layer_2_weights[12][0] = 0;
        layer_2_weights[13][0] = 0;
        layer_2_weights[14][0] = 1;
        layer_2_weights[15][0] = 5;
        layer_2_weights[0][1] = 7;
        layer_2_weights[1][1] = -3;
        layer_2_weights[2][1] = 5;
        layer_2_weights[3][1] = -5;
        layer_2_weights[4][1] = -4;
        layer_2_weights[5][1] = 3;
        layer_2_weights[6][1] = 4;
        layer_2_weights[7][1] = 3;
        layer_2_weights[8][1] = -5;
        layer_2_weights[9][1] = 2;
        layer_2_weights[10][1] = -3;
        layer_2_weights[11][1] = -10;
        layer_2_weights[12][1] = 1;
        layer_2_weights[13][1] = 4;
        layer_2_weights[14][1] = -1;
        layer_2_weights[15][1] = 5;
        layer_2_weights[0][2] = 0;
        layer_2_weights[1][2] = 0;
        layer_2_weights[2][2] = 0;
        layer_2_weights[3][2] = 0;
        layer_2_weights[4][2] = 3;
        layer_2_weights[5][2] = 2;
        layer_2_weights[6][2] = 3;
        layer_2_weights[7][2] = 3;
        layer_2_weights[8][2] = -2;
        layer_2_weights[9][2] = -1;
        layer_2_weights[10][2] = -3;
        layer_2_weights[11][2] = 2;
        layer_2_weights[12][2] = -3;
        layer_2_weights[13][2] = 8;
        layer_2_weights[14][2] = 4;
        layer_2_weights[15][2] = -11;
        layer_2_weights[0][3] = -4;
        layer_2_weights[1][3] = 4;
        layer_2_weights[2][3] = 2;
        layer_2_weights[3][3] = -8;
        layer_2_weights[4][3] = 3;
        layer_2_weights[5][3] = 2;
        layer_2_weights[6][3] = -1;
        layer_2_weights[7][3] = 4;
        layer_2_weights[8][3] = 3;
        layer_2_weights[9][3] = 3;
        layer_2_weights[10][3] = -1;
        layer_2_weights[11][3] = -1;
        layer_2_weights[12][3] = -4;
        layer_2_weights[13][3] = -2;
        layer_2_weights[14][3] = -3;
        layer_2_weights[15][3] = -5;
        layer_2_weights[0][4] = -3;
        layer_2_weights[1][4] = -7;
        layer_2_weights[2][4] = -15;
        layer_2_weights[3][4] = 3;
        layer_2_weights[4][4] = 2;
        layer_2_weights[5][4] = -4;
        layer_2_weights[6][4] = -3;
        layer_2_weights[7][4] = -12;
        layer_2_weights[8][4] = 2;
        layer_2_weights[9][4] = 4;
        layer_2_weights[10][4] = 3;
        layer_2_weights[11][4] = 1;
        layer_2_weights[12][4] = 1;
        layer_2_weights[13][4] = -9;
        layer_2_weights[14][4] = 0;
        layer_2_weights[15][4] = 5;
        layer_2_weights[0][5] = -5;
        layer_2_weights[1][5] = 2;
        layer_2_weights[2][5] = 6;
        layer_2_weights[3][5] = 3;
        layer_2_weights[4][5] = -8;
        layer_2_weights[5][5] = -3;
        layer_2_weights[6][5] = 5;
        layer_2_weights[7][5] = -3;
        layer_2_weights[8][5] = 4;
        layer_2_weights[9][5] = 2;
        layer_2_weights[10][5] = -2;
        layer_2_weights[11][5] = -2;
        layer_2_weights[12][5] = 3;
        layer_2_weights[13][5] = -5;
        layer_2_weights[14][5] = -3;
        layer_2_weights[15][5] = -3;
        layer_2_weights[0][6] = 6;
        layer_2_weights[1][6] = -4;
        layer_2_weights[2][6] = 0;
        layer_2_weights[3][6] = -1;
        layer_2_weights[4][6] = -3;
        layer_2_weights[5][6] = -3;
        layer_2_weights[6][6] = -4;
        layer_2_weights[7][6] = -5;
        layer_2_weights[8][6] = 4;
        layer_2_weights[9][6] = -4;
        layer_2_weights[10][6] = -3;
        layer_2_weights[11][6] = 4;
        layer_2_weights[12][6] = 6;
        layer_2_weights[13][6] = -1;
        layer_2_weights[14][6] = 2;
        layer_2_weights[15][6] = 2;
        layer_2_weights[0][7] = 1;
        layer_2_weights[1][7] = 3;
        layer_2_weights[2][7] = -1;
        layer_2_weights[3][7] = 5;
        layer_2_weights[4][7] = 3;
        layer_2_weights[5][7] = 4;
        layer_2_weights[6][7] = -3;
        layer_2_weights[7][7] = 0;
        layer_2_weights[8][7] = -5;
        layer_2_weights[9][7] = 0;
        layer_2_weights[10][7] = 4;
        layer_2_weights[11][7] = -1;
        layer_2_weights[12][7] = -5;
        layer_2_weights[13][7] = 3;
        layer_2_weights[14][7] = -6;
        layer_2_weights[15][7] = 3;
        layer_2_weights[0][8] = 0;
        layer_2_weights[1][8] = 2;
        layer_2_weights[2][8] = -6;
        layer_2_weights[3][8] = -1;
        layer_2_weights[4][8] = -1;
        layer_2_weights[5][8] = 1;
        layer_2_weights[6][8] = -2;
        layer_2_weights[7][8] = -5;
        layer_2_weights[8][8] = 1;
        layer_2_weights[9][8] = 1;
        layer_2_weights[10][8] = 2;
        layer_2_weights[11][8] = -6;
        layer_2_weights[12][8] = 4;
        layer_2_weights[13][8] = 3;
        layer_2_weights[14][8] = 3;
        layer_2_weights[15][8] = -4;
        layer_2_weights[0][9] = -7;
        layer_2_weights[1][9] = 3;
        layer_2_weights[2][9] = -5;
        layer_2_weights[3][9] = -4;
        layer_2_weights[4][9] = 6;
        layer_2_weights[5][9] = -12;
        layer_2_weights[6][9] = 1;
        layer_2_weights[7][9] = -4;
        layer_2_weights[8][9] = -4;
        layer_2_weights[9][9] = 2;
        layer_2_weights[10][9] = 4;
        layer_2_weights[11][9] = 4;
        layer_2_weights[12][9] = 3;
        layer_2_weights[13][9] = -6;
        layer_2_weights[14][9] = 0;
        layer_2_weights[15][9] = 1;
        layer_2_biases[0] = -6;
        layer_2_biases[1] = 2;
        layer_2_biases[2] = 0;
        layer_2_biases[3] = -2;
        layer_2_biases[4] = 2;
        layer_2_biases[5] = 7;
        layer_2_biases[6] = -1;
        layer_2_biases[7] = 1;
        layer_2_biases[8] = -4;
        layer_2_biases[9] = -1;
    end

    integer i, j, k;
    always @(*) begin
        if (predict) begin

            // Layer 1 Computation
            for (j = 0; j < 16; j = j + 1) begin
                layer_1_outputs[j] = layer_1_biases[j]; // Initialize with bias
                for (k = 0; k < 783; k = k + 1) begin
                    if (inp[k] == 1)
                        layer_1_outputs[j] = layer_1_outputs[j] + layer_1_weights[k][j];
                end
            end

            // Layer 2 Computation
            for (j = 0; j < 10; j = j + 1) begin
                layer_2_outputs[j] = layer_2_biases[j]; // Initialize with bias
                for (k = 0; k < 16; k = k + 1) begin
                    layer_2_outputs[j] = layer_2_outputs[j] + layer_1_outputs[k] * layer_2_weights[k][j];
                end
                // Apply ReLU
                if (layer_2_outputs[j] < 0)
                    layer_2_outputs[j] = 0;
            end

            // Winner-takes-all logic
            max_val = layer_2_outputs[0];
            max_idx = 0;
            for (i = 1; i < 10; i = i + 1) begin
                if (layer_2_outputs[i] > max_val) begin
                    max_val = layer_2_outputs[i];
                    max_idx = i;
                end
            end
            class = max_idx;

        end else begin
            class = 10;
        end
    end

endmodule
