module MLP_model (
    input predict,
    input [143:0] inp,
    output reg [3:0] class
);

    // Layer 1: Dense
    reg signed [7:0] layer_1_weights [143:0][15:0];
    reg signed [7:0] layer_1_biases [15:0];
    reg signed [8:0] layer_1_outputs [15:0];

    // Layer 2: Dense
    reg signed [7:0] layer_2_weights [15:0][9:0];
    reg signed [7:0] layer_2_biases [9:0];
    reg signed [17:0] layer_2_outputs [9:0];

    reg signed [17:0] max_val;
    reg [3:0] max_idx;

    initial begin
        layer_1_weights[0][0] = 2;
        layer_1_weights[1][0] = 2;
        layer_1_weights[2][0] = 1;
        layer_1_weights[3][0] = 11;
        layer_1_weights[4][0] = 18;
        layer_1_weights[5][0] = 4;
        layer_1_weights[6][0] = -11;
        layer_1_weights[7][0] = 8;
        layer_1_weights[8][0] = 2;
        layer_1_weights[9][0] = 16;
        layer_1_weights[10][0] = 2;
        layer_1_weights[11][0] = -2;
        layer_1_weights[12][0] = 2;
        layer_1_weights[13][0] = -2;
        layer_1_weights[14][0] = 4;
        layer_1_weights[15][0] = 2;
        layer_1_weights[16][0] = 11;
        layer_1_weights[17][0] = -2;
        layer_1_weights[18][0] = -6;
        layer_1_weights[19][0] = 0;
        layer_1_weights[20][0] = 0;
        layer_1_weights[21][0] = -5;
        layer_1_weights[22][0] = -1;
        layer_1_weights[23][0] = 6;
        layer_1_weights[24][0] = 1;
        layer_1_weights[25][0] = -3;
        layer_1_weights[26][0] = 1;
        layer_1_weights[27][0] = -1;
        layer_1_weights[28][0] = 2;
        layer_1_weights[29][0] = -3;
        layer_1_weights[30][0] = -2;
        layer_1_weights[31][0] = -5;
        layer_1_weights[32][0] = -5;
        layer_1_weights[33][0] = -5;
        layer_1_weights[34][0] = -3;
        layer_1_weights[35][0] = 10;
        layer_1_weights[36][0] = 1;
        layer_1_weights[37][0] = 2;
        layer_1_weights[38][0] = 1;
        layer_1_weights[39][0] = 1;
        layer_1_weights[40][0] = 2;
        layer_1_weights[41][0] = -1;
        layer_1_weights[42][0] = -4;
        layer_1_weights[43][0] = -4;
        layer_1_weights[44][0] = -4;
        layer_1_weights[45][0] = -3;
        layer_1_weights[46][0] = -3;
        layer_1_weights[47][0] = 7;
        layer_1_weights[48][0] = 1;
        layer_1_weights[49][0] = 3;
        layer_1_weights[50][0] = -2;
        layer_1_weights[51][0] = 0;
        layer_1_weights[52][0] = -6;
        layer_1_weights[53][0] = -2;
        layer_1_weights[54][0] = 0;
        layer_1_weights[55][0] = -3;
        layer_1_weights[56][0] = -5;
        layer_1_weights[57][0] = -2;
        layer_1_weights[58][0] = -12;
        layer_1_weights[59][0] = -11;
        layer_1_weights[60][0] = -4;
        layer_1_weights[61][0] = -16;
        layer_1_weights[62][0] = -8;
        layer_1_weights[63][0] = -9;
        layer_1_weights[64][0] = -1;
        layer_1_weights[65][0] = 5;
        layer_1_weights[66][0] = 4;
        layer_1_weights[67][0] = -3;
        layer_1_weights[68][0] = 0;
        layer_1_weights[69][0] = 1;
        layer_1_weights[70][0] = 4;
        layer_1_weights[71][0] = 9;
        layer_1_weights[72][0] = -4;
        layer_1_weights[73][0] = -12;
        layer_1_weights[74][0] = -4;
        layer_1_weights[75][0] = 2;
        layer_1_weights[76][0] = 9;
        layer_1_weights[77][0] = 15;
        layer_1_weights[78][0] = 11;
        layer_1_weights[79][0] = 3;
        layer_1_weights[80][0] = 7;
        layer_1_weights[81][0] = 12;
        layer_1_weights[82][0] = 12;
        layer_1_weights[83][0] = 23;
        layer_1_weights[84][0] = -9;
        layer_1_weights[85][0] = 5;
        layer_1_weights[86][0] = 9;
        layer_1_weights[87][0] = 9;
        layer_1_weights[88][0] = -3;
        layer_1_weights[89][0] = -1;
        layer_1_weights[90][0] = 8;
        layer_1_weights[91][0] = 10;
        layer_1_weights[92][0] = 11;
        layer_1_weights[93][0] = 11;
        layer_1_weights[94][0] = 12;
        layer_1_weights[95][0] = 10;
        layer_1_weights[96][0] = -6;
        layer_1_weights[97][0] = 1;
        layer_1_weights[98][0] = -5;
        layer_1_weights[99][0] = 5;
        layer_1_weights[100][0] = 0;
        layer_1_weights[101][0] = 0;
        layer_1_weights[102][0] = 3;
        layer_1_weights[103][0] = 4;
        layer_1_weights[104][0] = 1;
        layer_1_weights[105][0] = 5;
        layer_1_weights[106][0] = 2;
        layer_1_weights[107][0] = 7;
        layer_1_weights[108][0] = 8;
        layer_1_weights[109][0] = 0;
        layer_1_weights[110][0] = -5;
        layer_1_weights[111][0] = 1;
        layer_1_weights[112][0] = 1;
        layer_1_weights[113][0] = -3;
        layer_1_weights[114][0] = -9;
        layer_1_weights[115][0] = -7;
        layer_1_weights[116][0] = -14;
        layer_1_weights[117][0] = -12;
        layer_1_weights[118][0] = -11;
        layer_1_weights[119][0] = -6;
        layer_1_weights[120][0] = 1;
        layer_1_weights[121][0] = 0;
        layer_1_weights[122][0] = -8;
        layer_1_weights[123][0] = -8;
        layer_1_weights[124][0] = -4;
        layer_1_weights[125][0] = -8;
        layer_1_weights[126][0] = -7;
        layer_1_weights[127][0] = -12;
        layer_1_weights[128][0] = -16;
        layer_1_weights[129][0] = -4;
        layer_1_weights[130][0] = -22;
        layer_1_weights[131][0] = 13;
        layer_1_weights[132][0] = 3;
        layer_1_weights[133][0] = -2;
        layer_1_weights[134][0] = -19;
        layer_1_weights[135][0] = -25;
        layer_1_weights[136][0] = -16;
        layer_1_weights[137][0] = -14;
        layer_1_weights[138][0] = -16;
        layer_1_weights[139][0] = -11;
        layer_1_weights[140][0] = -3;
        layer_1_weights[141][0] = -8;
        layer_1_weights[142][0] = 0;
        layer_1_weights[143][0] = 3;
        layer_1_weights[0][1] = -3;
        layer_1_weights[1][1] = -3;
        layer_1_weights[2][1] = 7;
        layer_1_weights[3][1] = 12;
        layer_1_weights[4][1] = 17;
        layer_1_weights[5][1] = 1;
        layer_1_weights[6][1] = -7;
        layer_1_weights[7][1] = 9;
        layer_1_weights[8][1] = 0;
        layer_1_weights[9][1] = 22;
        layer_1_weights[10][1] = 0;
        layer_1_weights[11][1] = 2;
        layer_1_weights[12][1] = 2;
        layer_1_weights[13][1] = 3;
        layer_1_weights[14][1] = -5;
        layer_1_weights[15][1] = -2;
        layer_1_weights[16][1] = 3;
        layer_1_weights[17][1] = 4;
        layer_1_weights[18][1] = 7;
        layer_1_weights[19][1] = 5;
        layer_1_weights[20][1] = 3;
        layer_1_weights[21][1] = -3;
        layer_1_weights[22][1] = 11;
        layer_1_weights[23][1] = 8;
        layer_1_weights[24][1] = 0;
        layer_1_weights[25][1] = 6;
        layer_1_weights[26][1] = -8;
        layer_1_weights[27][1] = 4;
        layer_1_weights[28][1] = -5;
        layer_1_weights[29][1] = -1;
        layer_1_weights[30][1] = 1;
        layer_1_weights[31][1] = 0;
        layer_1_weights[32][1] = -2;
        layer_1_weights[33][1] = 2;
        layer_1_weights[34][1] = 6;
        layer_1_weights[35][1] = 12;
        layer_1_weights[36][1] = -14;
        layer_1_weights[37][1] = 1;
        layer_1_weights[38][1] = -5;
        layer_1_weights[39][1] = -2;
        layer_1_weights[40][1] = -2;
        layer_1_weights[41][1] = -1;
        layer_1_weights[42][1] = 2;
        layer_1_weights[43][1] = 2;
        layer_1_weights[44][1] = -1;
        layer_1_weights[45][1] = -2;
        layer_1_weights[46][1] = -1;
        layer_1_weights[47][1] = 12;
        layer_1_weights[48][1] = -20;
        layer_1_weights[49][1] = -5;
        layer_1_weights[50][1] = 0;
        layer_1_weights[51][1] = 0;
        layer_1_weights[52][1] = -1;
        layer_1_weights[53][1] = -14;
        layer_1_weights[54][1] = -12;
        layer_1_weights[55][1] = -3;
        layer_1_weights[56][1] = -1;
        layer_1_weights[57][1] = 1;
        layer_1_weights[58][1] = -9;
        layer_1_weights[59][1] = -10;
        layer_1_weights[60][1] = -10;
        layer_1_weights[61][1] = 0;
        layer_1_weights[62][1] = 5;
        layer_1_weights[63][1] = 10;
        layer_1_weights[64][1] = 8;
        layer_1_weights[65][1] = -8;
        layer_1_weights[66][1] = -6;
        layer_1_weights[67][1] = 4;
        layer_1_weights[68][1] = 5;
        layer_1_weights[69][1] = 2;
        layer_1_weights[70][1] = 4;
        layer_1_weights[71][1] = -8;
        layer_1_weights[72][1] = 2;
        layer_1_weights[73][1] = -4;
        layer_1_weights[74][1] = 3;
        layer_1_weights[75][1] = 6;
        layer_1_weights[76][1] = 11;
        layer_1_weights[77][1] = 17;
        layer_1_weights[78][1] = 4;
        layer_1_weights[79][1] = 4;
        layer_1_weights[80][1] = 2;
        layer_1_weights[81][1] = -4;
        layer_1_weights[82][1] = 1;
        layer_1_weights[83][1] = 10;
        layer_1_weights[84][1] = -3;
        layer_1_weights[85][1] = -1;
        layer_1_weights[86][1] = 6;
        layer_1_weights[87][1] = 0;
        layer_1_weights[88][1] = 7;
        layer_1_weights[89][1] = 16;
        layer_1_weights[90][1] = 4;
        layer_1_weights[91][1] = 3;
        layer_1_weights[92][1] = 0;
        layer_1_weights[93][1] = -6;
        layer_1_weights[94][1] = 0;
        layer_1_weights[95][1] = -9;
        layer_1_weights[96][1] = 11;
        layer_1_weights[97][1] = -4;
        layer_1_weights[98][1] = -2;
        layer_1_weights[99][1] = -5;
        layer_1_weights[100][1] = 5;
        layer_1_weights[101][1] = 5;
        layer_1_weights[102][1] = 4;
        layer_1_weights[103][1] = 10;
        layer_1_weights[104][1] = 5;
        layer_1_weights[105][1] = 7;
        layer_1_weights[106][1] = -5;
        layer_1_weights[107][1] = 5;
        layer_1_weights[108][1] = 12;
        layer_1_weights[109][1] = -2;
        layer_1_weights[110][1] = -16;
        layer_1_weights[111][1] = -8;
        layer_1_weights[112][1] = -5;
        layer_1_weights[113][1] = -1;
        layer_1_weights[114][1] = 3;
        layer_1_weights[115][1] = 4;
        layer_1_weights[116][1] = 9;
        layer_1_weights[117][1] = 1;
        layer_1_weights[118][1] = 13;
        layer_1_weights[119][1] = 0;
        layer_1_weights[120][1] = -3;
        layer_1_weights[121][1] = 12;
        layer_1_weights[122][1] = -6;
        layer_1_weights[123][1] = -12;
        layer_1_weights[124][1] = -8;
        layer_1_weights[125][1] = -8;
        layer_1_weights[126][1] = -5;
        layer_1_weights[127][1] = -1;
        layer_1_weights[128][1] = 6;
        layer_1_weights[129][1] = 16;
        layer_1_weights[130][1] = 10;
        layer_1_weights[131][1] = -10;
        layer_1_weights[132][1] = -3;
        layer_1_weights[133][1] = 1;
        layer_1_weights[134][1] = 10;
        layer_1_weights[135][1] = 5;
        layer_1_weights[136][1] = 6;
        layer_1_weights[137][1] = 3;
        layer_1_weights[138][1] = -1;
        layer_1_weights[139][1] = -4;
        layer_1_weights[140][1] = -6;
        layer_1_weights[141][1] = -3;
        layer_1_weights[142][1] = 1;
        layer_1_weights[143][1] = -1;
        layer_1_weights[0][2] = 3;
        layer_1_weights[1][2] = 1;
        layer_1_weights[2][2] = 2;
        layer_1_weights[3][2] = 3;
        layer_1_weights[4][2] = -12;
        layer_1_weights[5][2] = 3;
        layer_1_weights[6][2] = 9;
        layer_1_weights[7][2] = 5;
        layer_1_weights[8][2] = 8;
        layer_1_weights[9][2] = 12;
        layer_1_weights[10][2] = -1;
        layer_1_weights[11][2] = -1;
        layer_1_weights[12][2] = -3;
        layer_1_weights[13][2] = 3;
        layer_1_weights[14][2] = 5;
        layer_1_weights[15][2] = -2;
        layer_1_weights[16][2] = 3;
        layer_1_weights[17][2] = 1;
        layer_1_weights[18][2] = 2;
        layer_1_weights[19][2] = -2;
        layer_1_weights[20][2] = -3;
        layer_1_weights[21][2] = -11;
        layer_1_weights[22][2] = -16;
        layer_1_weights[23][2] = 10;
        layer_1_weights[24][2] = 2;
        layer_1_weights[25][2] = 9;
        layer_1_weights[26][2] = -9;
        layer_1_weights[27][2] = -4;
        layer_1_weights[28][2] = -2;
        layer_1_weights[29][2] = -2;
        layer_1_weights[30][2] = 0;
        layer_1_weights[31][2] = 0;
        layer_1_weights[32][2] = -3;
        layer_1_weights[33][2] = -6;
        layer_1_weights[34][2] = -10;
        layer_1_weights[35][2] = 5;
        layer_1_weights[36][2] = -8;
        layer_1_weights[37][2] = 2;
        layer_1_weights[38][2] = 4;
        layer_1_weights[39][2] = 5;
        layer_1_weights[40][2] = 1;
        layer_1_weights[41][2] = 1;
        layer_1_weights[42][2] = 11;
        layer_1_weights[43][2] = 6;
        layer_1_weights[44][2] = -1;
        layer_1_weights[45][2] = -2;
        layer_1_weights[46][2] = -6;
        layer_1_weights[47][2] = -7;
        layer_1_weights[48][2] = -1;
        layer_1_weights[49][2] = 4;
        layer_1_weights[50][2] = 5;
        layer_1_weights[51][2] = 3;
        layer_1_weights[52][2] = -7;
        layer_1_weights[53][2] = 1;
        layer_1_weights[54][2] = 8;
        layer_1_weights[55][2] = 1;
        layer_1_weights[56][2] = 6;
        layer_1_weights[57][2] = 5;
        layer_1_weights[58][2] = 2;
        layer_1_weights[59][2] = -5;
        layer_1_weights[60][2] = -17;
        layer_1_weights[61][2] = 2;
        layer_1_weights[62][2] = 2;
        layer_1_weights[63][2] = 1;
        layer_1_weights[64][2] = -4;
        layer_1_weights[65][2] = 3;
        layer_1_weights[66][2] = 14;
        layer_1_weights[67][2] = 0;
        layer_1_weights[68][2] = 3;
        layer_1_weights[69][2] = -3;
        layer_1_weights[70][2] = -4;
        layer_1_weights[71][2] = 10;
        layer_1_weights[72][2] = 5;
        layer_1_weights[73][2] = -3;
        layer_1_weights[74][2] = -6;
        layer_1_weights[75][2] = -3;
        layer_1_weights[76][2] = 5;
        layer_1_weights[77][2] = 17;
        layer_1_weights[78][2] = 9;
        layer_1_weights[79][2] = 0;
        layer_1_weights[80][2] = -3;
        layer_1_weights[81][2] = -1;
        layer_1_weights[82][2] = -3;
        layer_1_weights[83][2] = -8;
        layer_1_weights[84][2] = 22;
        layer_1_weights[85][2] = 3;
        layer_1_weights[86][2] = -5;
        layer_1_weights[87][2] = 0;
        layer_1_weights[88][2] = 15;
        layer_1_weights[89][2] = 10;
        layer_1_weights[90][2] = 0;
        layer_1_weights[91][2] = -2;
        layer_1_weights[92][2] = -2;
        layer_1_weights[93][2] = 0;
        layer_1_weights[94][2] = 2;
        layer_1_weights[95][2] = -11;
        layer_1_weights[96][2] = -4;
        layer_1_weights[97][2] = -4;
        layer_1_weights[98][2] = -1;
        layer_1_weights[99][2] = -1;
        layer_1_weights[100][2] = -1;
        layer_1_weights[101][2] = -7;
        layer_1_weights[102][2] = -6;
        layer_1_weights[103][2] = 3;
        layer_1_weights[104][2] = 3;
        layer_1_weights[105][2] = 5;
        layer_1_weights[106][2] = 5;
        layer_1_weights[107][2] = -3;
        layer_1_weights[108][2] = 8;
        layer_1_weights[109][2] = 1;
        layer_1_weights[110][2] = 5;
        layer_1_weights[111][2] = 3;
        layer_1_weights[112][2] = -1;
        layer_1_weights[113][2] = 2;
        layer_1_weights[114][2] = 2;
        layer_1_weights[115][2] = 1;
        layer_1_weights[116][2] = -1;
        layer_1_weights[117][2] = -4;
        layer_1_weights[118][2] = -1;
        layer_1_weights[119][2] = -10;
        layer_1_weights[120][2] = -3;
        layer_1_weights[121][2] = -1;
        layer_1_weights[122][2] = 2;
        layer_1_weights[123][2] = 5;
        layer_1_weights[124][2] = 7;
        layer_1_weights[125][2] = 7;
        layer_1_weights[126][2] = 2;
        layer_1_weights[127][2] = -3;
        layer_1_weights[128][2] = -3;
        layer_1_weights[129][2] = -2;
        layer_1_weights[130][2] = -7;
        layer_1_weights[131][2] = -14;
        layer_1_weights[132][2] = -2;
        layer_1_weights[133][2] = -1;
        layer_1_weights[134][2] = -1;
        layer_1_weights[135][2] = 5;
        layer_1_weights[136][2] = 5;
        layer_1_weights[137][2] = 6;
        layer_1_weights[138][2] = -1;
        layer_1_weights[139][2] = 5;
        layer_1_weights[140][2] = 8;
        layer_1_weights[141][2] = -2;
        layer_1_weights[142][2] = 3;
        layer_1_weights[143][2] = 0;
        layer_1_weights[0][3] = 1;
        layer_1_weights[1][3] = 0;
        layer_1_weights[2][3] = 4;
        layer_1_weights[3][3] = -1;
        layer_1_weights[4][3] = -10;
        layer_1_weights[5][3] = -1;
        layer_1_weights[6][3] = 20;
        layer_1_weights[7][3] = 14;
        layer_1_weights[8][3] = 17;
        layer_1_weights[9][3] = -10;
        layer_1_weights[10][3] = -3;
        layer_1_weights[11][3] = 1;
        layer_1_weights[12][3] = 3;
        layer_1_weights[13][3] = 0;
        layer_1_weights[14][3] = -1;
        layer_1_weights[15][3] = -6;
        layer_1_weights[16][3] = -3;
        layer_1_weights[17][3] = 1;
        layer_1_weights[18][3] = 3;
        layer_1_weights[19][3] = 5;
        layer_1_weights[20][3] = 8;
        layer_1_weights[21][3] = 9;
        layer_1_weights[22][3] = 0;
        layer_1_weights[23][3] = 5;
        layer_1_weights[24][3] = -3;
        layer_1_weights[25][3] = 1;
        layer_1_weights[26][3] = 1;
        layer_1_weights[27][3] = 2;
        layer_1_weights[28][3] = 1;
        layer_1_weights[29][3] = 2;
        layer_1_weights[30][3] = 3;
        layer_1_weights[31][3] = 5;
        layer_1_weights[32][3] = 6;
        layer_1_weights[33][3] = 5;
        layer_1_weights[34][3] = 7;
        layer_1_weights[35][3] = 1;
        layer_1_weights[36][3] = -2;
        layer_1_weights[37][3] = -1;
        layer_1_weights[38][3] = 0;
        layer_1_weights[39][3] = 0;
        layer_1_weights[40][3] = 2;
        layer_1_weights[41][3] = 11;
        layer_1_weights[42][3] = 12;
        layer_1_weights[43][3] = 1;
        layer_1_weights[44][3] = 1;
        layer_1_weights[45][3] = 4;
        layer_1_weights[46][3] = 8;
        layer_1_weights[47][3] = 9;
        layer_1_weights[48][3] = 4;
        layer_1_weights[49][3] = 0;
        layer_1_weights[50][3] = -1;
        layer_1_weights[51][3] = 1;
        layer_1_weights[52][3] = 0;
        layer_1_weights[53][3] = 4;
        layer_1_weights[54][3] = -6;
        layer_1_weights[55][3] = -13;
        layer_1_weights[56][3] = -13;
        layer_1_weights[57][3] = -19;
        layer_1_weights[58][3] = -10;
        layer_1_weights[59][3] = 9;
        layer_1_weights[60][3] = -16;
        layer_1_weights[61][3] = 2;
        layer_1_weights[62][3] = -2;
        layer_1_weights[63][3] = 1;
        layer_1_weights[64][3] = 1;
        layer_1_weights[65][3] = 2;
        layer_1_weights[66][3] = -3;
        layer_1_weights[67][3] = -10;
        layer_1_weights[68][3] = -1;
        layer_1_weights[69][3] = -11;
        layer_1_weights[70][3] = -9;
        layer_1_weights[71][3] = -16;
        layer_1_weights[72][3] = -6;
        layer_1_weights[73][3] = 1;
        layer_1_weights[74][3] = -2;
        layer_1_weights[75][3] = 3;
        layer_1_weights[76][3] = 3;
        layer_1_weights[77][3] = -1;
        layer_1_weights[78][3] = -4;
        layer_1_weights[79][3] = -4;
        layer_1_weights[80][3] = -2;
        layer_1_weights[81][3] = -2;
        layer_1_weights[82][3] = 1;
        layer_1_weights[83][3] = -24;
        layer_1_weights[84][3] = 4;
        layer_1_weights[85][3] = 1;
        layer_1_weights[86][3] = -9;
        layer_1_weights[87][3] = -8;
        layer_1_weights[88][3] = -7;
        layer_1_weights[89][3] = -2;
        layer_1_weights[90][3] = -4;
        layer_1_weights[91][3] = -3;
        layer_1_weights[92][3] = -3;
        layer_1_weights[93][3] = -2;
        layer_1_weights[94][3] = -2;
        layer_1_weights[95][3] = -11;
        layer_1_weights[96][3] = -2;
        layer_1_weights[97][3] = 1;
        layer_1_weights[98][3] = 7;
        layer_1_weights[99][3] = -4;
        layer_1_weights[100][3] = -10;
        layer_1_weights[101][3] = -3;
        layer_1_weights[102][3] = 3;
        layer_1_weights[103][3] = 9;
        layer_1_weights[104][3] = 5;
        layer_1_weights[105][3] = 9;
        layer_1_weights[106][3] = 5;
        layer_1_weights[107][3] = 5;
        layer_1_weights[108][3] = 5;
        layer_1_weights[109][3] = 11;
        layer_1_weights[110][3] = 9;
        layer_1_weights[111][3] = 9;
        layer_1_weights[112][3] = 9;
        layer_1_weights[113][3] = 5;
        layer_1_weights[114][3] = 8;
        layer_1_weights[115][3] = 9;
        layer_1_weights[116][3] = 12;
        layer_1_weights[117][3] = 14;
        layer_1_weights[118][3] = 17;
        layer_1_weights[119][3] = 17;
        layer_1_weights[120][3] = -1;
        layer_1_weights[121][3] = 15;
        layer_1_weights[122][3] = 8;
        layer_1_weights[123][3] = 7;
        layer_1_weights[124][3] = 9;
        layer_1_weights[125][3] = 6;
        layer_1_weights[126][3] = 6;
        layer_1_weights[127][3] = 4;
        layer_1_weights[128][3] = 3;
        layer_1_weights[129][3] = 2;
        layer_1_weights[130][3] = 11;
        layer_1_weights[131][3] = 6;
        layer_1_weights[132][3] = 1;
        layer_1_weights[133][3] = 0;
        layer_1_weights[134][3] = 8;
        layer_1_weights[135][3] = 2;
        layer_1_weights[136][3] = 2;
        layer_1_weights[137][3] = -4;
        layer_1_weights[138][3] = 1;
        layer_1_weights[139][3] = -3;
        layer_1_weights[140][3] = -6;
        layer_1_weights[141][3] = 5;
        layer_1_weights[142][3] = -1;
        layer_1_weights[143][3] = 0;
        layer_1_weights[0][4] = -2;
        layer_1_weights[1][4] = 0;
        layer_1_weights[2][4] = 7;
        layer_1_weights[3][4] = 14;
        layer_1_weights[4][4] = 27;
        layer_1_weights[5][4] = -2;
        layer_1_weights[6][4] = -2;
        layer_1_weights[7][4] = -8;
        layer_1_weights[8][4] = -3;
        layer_1_weights[9][4] = -7;
        layer_1_weights[10][4] = -1;
        layer_1_weights[11][4] = 1;
        layer_1_weights[12][4] = 2;
        layer_1_weights[13][4] = 2;
        layer_1_weights[14][4] = -15;
        layer_1_weights[15][4] = -10;
        layer_1_weights[16][4] = -8;
        layer_1_weights[17][4] = -7;
        layer_1_weights[18][4] = -4;
        layer_1_weights[19][4] = 3;
        layer_1_weights[20][4] = 11;
        layer_1_weights[21][4] = 15;
        layer_1_weights[22][4] = 15;
        layer_1_weights[23][4] = -5;
        layer_1_weights[24][4] = 3;
        layer_1_weights[25][4] = -8;
        layer_1_weights[26][4] = -1;
        layer_1_weights[27][4] = 1;
        layer_1_weights[28][4] = 1;
        layer_1_weights[29][4] = 2;
        layer_1_weights[30][4] = 2;
        layer_1_weights[31][4] = 2;
        layer_1_weights[32][4] = 5;
        layer_1_weights[33][4] = 11;
        layer_1_weights[34][4] = 16;
        layer_1_weights[35][4] = 15;
        layer_1_weights[36][4] = -8;
        layer_1_weights[37][4] = -6;
        layer_1_weights[38][4] = 1;
        layer_1_weights[39][4] = 0;
        layer_1_weights[40][4] = 5;
        layer_1_weights[41][4] = 2;
        layer_1_weights[42][4] = -12;
        layer_1_weights[43][4] = -5;
        layer_1_weights[44][4] = 4;
        layer_1_weights[45][4] = 8;
        layer_1_weights[46][4] = 18;
        layer_1_weights[47][4] = 27;
        layer_1_weights[48][4] = -10;
        layer_1_weights[49][4] = 2;
        layer_1_weights[50][4] = -7;
        layer_1_weights[51][4] = 0;
        layer_1_weights[52][4] = 5;
        layer_1_weights[53][4] = 1;
        layer_1_weights[54][4] = -12;
        layer_1_weights[55][4] = -7;
        layer_1_weights[56][4] = -8;
        layer_1_weights[57][4] = -8;
        layer_1_weights[58][4] = 5;
        layer_1_weights[59][4] = 8;
        layer_1_weights[60][4] = -4;
        layer_1_weights[61][4] = -5;
        layer_1_weights[62][4] = 2;
        layer_1_weights[63][4] = 2;
        layer_1_weights[64][4] = 8;
        layer_1_weights[65][4] = 10;
        layer_1_weights[66][4] = 3;
        layer_1_weights[67][4] = 5;
        layer_1_weights[68][4] = -2;
        layer_1_weights[69][4] = 0;
        layer_1_weights[70][4] = 1;
        layer_1_weights[71][4] = -10;
        layer_1_weights[72][4] = 2;
        layer_1_weights[73][4] = -7;
        layer_1_weights[74][4] = 5;
        layer_1_weights[75][4] = 7;
        layer_1_weights[76][4] = 9;
        layer_1_weights[77][4] = 7;
        layer_1_weights[78][4] = 12;
        layer_1_weights[79][4] = 8;
        layer_1_weights[80][4] = 0;
        layer_1_weights[81][4] = 4;
        layer_1_weights[82][4] = 6;
        layer_1_weights[83][4] = -4;
        layer_1_weights[84][4] = -12;
        layer_1_weights[85][4] = -6;
        layer_1_weights[86][4] = 2;
        layer_1_weights[87][4] = -2;
        layer_1_weights[88][4] = 4;
        layer_1_weights[89][4] = 5;
        layer_1_weights[90][4] = 8;
        layer_1_weights[91][4] = 0;
        layer_1_weights[92][4] = -5;
        layer_1_weights[93][4] = 2;
        layer_1_weights[94][4] = -4;
        layer_1_weights[95][4] = -4;
        layer_1_weights[96][4] = -10;
        layer_1_weights[97][4] = -7;
        layer_1_weights[98][4] = -6;
        layer_1_weights[99][4] = 1;
        layer_1_weights[100][4] = -3;
        layer_1_weights[101][4] = -3;
        layer_1_weights[102][4] = -1;
        layer_1_weights[103][4] = -6;
        layer_1_weights[104][4] = -5;
        layer_1_weights[105][4] = -9;
        layer_1_weights[106][4] = -4;
        layer_1_weights[107][4] = -4;
        layer_1_weights[108][4] = -3;
        layer_1_weights[109][4] = -1;
        layer_1_weights[110][4] = -10;
        layer_1_weights[111][4] = -3;
        layer_1_weights[112][4] = 3;
        layer_1_weights[113][4] = 5;
        layer_1_weights[114][4] = 1;
        layer_1_weights[115][4] = 1;
        layer_1_weights[116][4] = 2;
        layer_1_weights[117][4] = 8;
        layer_1_weights[118][4] = 1;
        layer_1_weights[119][4] = 12;
        layer_1_weights[120][4] = -2;
        layer_1_weights[121][4] = -11;
        layer_1_weights[122][4] = -2;
        layer_1_weights[123][4] = -1;
        layer_1_weights[124][4] = 0;
        layer_1_weights[125][4] = 3;
        layer_1_weights[126][4] = 6;
        layer_1_weights[127][4] = 6;
        layer_1_weights[128][4] = 3;
        layer_1_weights[129][4] = 1;
        layer_1_weights[130][4] = -3;
        layer_1_weights[131][4] = -12;
        layer_1_weights[132][4] = 0;
        layer_1_weights[133][4] = -4;
        layer_1_weights[134][4] = -34;
        layer_1_weights[135][4] = -5;
        layer_1_weights[136][4] = -8;
        layer_1_weights[137][4] = -9;
        layer_1_weights[138][4] = -9;
        layer_1_weights[139][4] = -11;
        layer_1_weights[140][4] = -13;
        layer_1_weights[141][4] = -5;
        layer_1_weights[142][4] = 2;
        layer_1_weights[143][4] = 1;
        layer_1_weights[0][5] = -2;
        layer_1_weights[1][5] = 0;
        layer_1_weights[2][5] = 1;
        layer_1_weights[3][5] = 0;
        layer_1_weights[4][5] = 1;
        layer_1_weights[5][5] = 0;
        layer_1_weights[6][5] = -14;
        layer_1_weights[7][5] = -13;
        layer_1_weights[8][5] = 8;
        layer_1_weights[9][5] = -1;
        layer_1_weights[10][5] = 3;
        layer_1_weights[11][5] = 2;
        layer_1_weights[12][5] = 1;
        layer_1_weights[13][5] = -1;
        layer_1_weights[14][5] = 7;
        layer_1_weights[15][5] = -8;
        layer_1_weights[16][5] = -7;
        layer_1_weights[17][5] = -11;
        layer_1_weights[18][5] = -6;
        layer_1_weights[19][5] = -3;
        layer_1_weights[20][5] = -22;
        layer_1_weights[21][5] = -13;
        layer_1_weights[22][5] = -16;
        layer_1_weights[23][5] = 2;
        layer_1_weights[24][5] = 2;
        layer_1_weights[25][5] = 2;
        layer_1_weights[26][5] = 1;
        layer_1_weights[27][5] = -3;
        layer_1_weights[28][5] = -2;
        layer_1_weights[29][5] = -2;
        layer_1_weights[30][5] = -8;
        layer_1_weights[31][5] = -8;
        layer_1_weights[32][5] = -5;
        layer_1_weights[33][5] = -5;
        layer_1_weights[34][5] = -4;
        layer_1_weights[35][5] = 1;
        layer_1_weights[36][5] = 8;
        layer_1_weights[37][5] = 1;
        layer_1_weights[38][5] = -2;
        layer_1_weights[39][5] = -3;
        layer_1_weights[40][5] = -8;
        layer_1_weights[41][5] = -5;
        layer_1_weights[42][5] = 4;
        layer_1_weights[43][5] = 12;
        layer_1_weights[44][5] = 10;
        layer_1_weights[45][5] = 12;
        layer_1_weights[46][5] = 9;
        layer_1_weights[47][5] = -2;
        layer_1_weights[48][5] = 3;
        layer_1_weights[49][5] = 0;
        layer_1_weights[50][5] = -4;
        layer_1_weights[51][5] = -4;
        layer_1_weights[52][5] = -3;
        layer_1_weights[53][5] = 3;
        layer_1_weights[54][5] = 8;
        layer_1_weights[55][5] = 10;
        layer_1_weights[56][5] = 11;
        layer_1_weights[57][5] = 13;
        layer_1_weights[58][5] = 13;
        layer_1_weights[59][5] = 10;
        layer_1_weights[60][5] = 14;
        layer_1_weights[61][5] = -3;
        layer_1_weights[62][5] = -6;
        layer_1_weights[63][5] = 3;
        layer_1_weights[64][5] = 6;
        layer_1_weights[65][5] = -1;
        layer_1_weights[66][5] = -4;
        layer_1_weights[67][5] = -10;
        layer_1_weights[68][5] = -16;
        layer_1_weights[69][5] = -14;
        layer_1_weights[70][5] = -8;
        layer_1_weights[71][5] = 23;
        layer_1_weights[72][5] = 4;
        layer_1_weights[73][5] = 0;
        layer_1_weights[74][5] = 5;
        layer_1_weights[75][5] = -1;
        layer_1_weights[76][5] = -1;
        layer_1_weights[77][5] = 6;
        layer_1_weights[78][5] = -5;
        layer_1_weights[79][5] = -3;
        layer_1_weights[80][5] = -8;
        layer_1_weights[81][5] = -16;
        layer_1_weights[82][5] = -6;
        layer_1_weights[83][5] = 5;
        layer_1_weights[84][5] = -1;
        layer_1_weights[85][5] = -5;
        layer_1_weights[86][5] = 5;
        layer_1_weights[87][5] = 0;
        layer_1_weights[88][5] = 1;
        layer_1_weights[89][5] = -3;
        layer_1_weights[90][5] = 0;
        layer_1_weights[91][5] = 2;
        layer_1_weights[92][5] = -3;
        layer_1_weights[93][5] = -7;
        layer_1_weights[94][5] = -6;
        layer_1_weights[95][5] = 12;
        layer_1_weights[96][5] = 7;
        layer_1_weights[97][5] = -10;
        layer_1_weights[98][5] = 2;
        layer_1_weights[99][5] = 3;
        layer_1_weights[100][5] = 0;
        layer_1_weights[101][5] = 3;
        layer_1_weights[102][5] = 2;
        layer_1_weights[103][5] = -3;
        layer_1_weights[104][5] = 0;
        layer_1_weights[105][5] = 1;
        layer_1_weights[106][5] = -16;
        layer_1_weights[107][5] = 7;
        layer_1_weights[108][5] = -2;
        layer_1_weights[109][5] = -10;
        layer_1_weights[110][5] = 1;
        layer_1_weights[111][5] = 1;
        layer_1_weights[112][5] = -1;
        layer_1_weights[113][5] = 0;
        layer_1_weights[114][5] = -5;
        layer_1_weights[115][5] = -3;
        layer_1_weights[116][5] = 0;
        layer_1_weights[117][5] = -5;
        layer_1_weights[118][5] = -9;
        layer_1_weights[119][5] = -13;
        layer_1_weights[120][5] = 2;
        layer_1_weights[121][5] = -8;
        layer_1_weights[122][5] = -6;
        layer_1_weights[123][5] = 1;
        layer_1_weights[124][5] = 4;
        layer_1_weights[125][5] = 1;
        layer_1_weights[126][5] = -1;
        layer_1_weights[127][5] = -2;
        layer_1_weights[128][5] = 2;
        layer_1_weights[129][5] = -5;
        layer_1_weights[130][5] = -12;
        layer_1_weights[131][5] = 1;
        layer_1_weights[132][5] = 1;
        layer_1_weights[133][5] = 9;
        layer_1_weights[134][5] = -3;
        layer_1_weights[135][5] = -8;
        layer_1_weights[136][5] = -3;
        layer_1_weights[137][5] = 4;
        layer_1_weights[138][5] = 1;
        layer_1_weights[139][5] = 4;
        layer_1_weights[140][5] = 8;
        layer_1_weights[141][5] = -12;
        layer_1_weights[142][5] = 2;
        layer_1_weights[143][5] = -2;
        layer_1_weights[0][6] = -2;
        layer_1_weights[1][6] = 2;
        layer_1_weights[2][6] = -9;
        layer_1_weights[3][6] = -18;
        layer_1_weights[4][6] = -33;
        layer_1_weights[5][6] = -13;
        layer_1_weights[6][6] = -11;
        layer_1_weights[7][6] = -4;
        layer_1_weights[8][6] = -29;
        layer_1_weights[9][6] = -18;
        layer_1_weights[10][6] = -3;
        layer_1_weights[11][6] = 1;
        layer_1_weights[12][6] = 1;
        layer_1_weights[13][6] = 0;
        layer_1_weights[14][6] = -10;
        layer_1_weights[15][6] = -30;
        layer_1_weights[16][6] = -33;
        layer_1_weights[17][6] = -31;
        layer_1_weights[18][6] = -22;
        layer_1_weights[19][6] = -15;
        layer_1_weights[20][6] = -8;
        layer_1_weights[21][6] = -9;
        layer_1_weights[22][6] = 2;
        layer_1_weights[23][6] = -2;
        layer_1_weights[24][6] = 3;
        layer_1_weights[25][6] = 1;
        layer_1_weights[26][6] = -7;
        layer_1_weights[27][6] = -1;
        layer_1_weights[28][6] = 0;
        layer_1_weights[29][6] = -5;
        layer_1_weights[30][6] = -4;
        layer_1_weights[31][6] = -1;
        layer_1_weights[32][6] = -1;
        layer_1_weights[33][6] = 4;
        layer_1_weights[34][6] = -3;
        layer_1_weights[35][6] = 6;
        layer_1_weights[36][6] = 10;
        layer_1_weights[37][6] = -8;
        layer_1_weights[38][6] = 6;
        layer_1_weights[39][6] = 9;
        layer_1_weights[40][6] = 10;
        layer_1_weights[41][6] = 10;
        layer_1_weights[42][6] = 8;
        layer_1_weights[43][6] = 4;
        layer_1_weights[44][6] = 2;
        layer_1_weights[45][6] = 5;
        layer_1_weights[46][6] = 7;
        layer_1_weights[47][6] = -1;
        layer_1_weights[48][6] = 8;
        layer_1_weights[49][6] = 3;
        layer_1_weights[50][6] = 7;
        layer_1_weights[51][6] = 13;
        layer_1_weights[52][6] = 5;
        layer_1_weights[53][6] = 6;
        layer_1_weights[54][6] = -2;
        layer_1_weights[55][6] = 1;
        layer_1_weights[56][6] = -1;
        layer_1_weights[57][6] = -1;
        layer_1_weights[58][6] = -6;
        layer_1_weights[59][6] = -6;
        layer_1_weights[60][6] = 15;
        layer_1_weights[61][6] = 6;
        layer_1_weights[62][6] = 6;
        layer_1_weights[63][6] = 9;
        layer_1_weights[64][6] = 1;
        layer_1_weights[65][6] = -4;
        layer_1_weights[66][6] = 1;
        layer_1_weights[67][6] = 3;
        layer_1_weights[68][6] = 5;
        layer_1_weights[69][6] = -1;
        layer_1_weights[70][6] = -5;
        layer_1_weights[71][6] = 6;
        layer_1_weights[72][6] = 3;
        layer_1_weights[73][6] = -1;
        layer_1_weights[74][6] = -3;
        layer_1_weights[75][6] = 6;
        layer_1_weights[76][6] = 5;
        layer_1_weights[77][6] = 3;
        layer_1_weights[78][6] = 5;
        layer_1_weights[79][6] = 8;
        layer_1_weights[80][6] = 9;
        layer_1_weights[81][6] = 4;
        layer_1_weights[82][6] = 5;
        layer_1_weights[83][6] = 8;
        layer_1_weights[84][6] = 5;
        layer_1_weights[85][6] = -1;
        layer_1_weights[86][6] = 4;
        layer_1_weights[87][6] = 0;
        layer_1_weights[88][6] = 0;
        layer_1_weights[89][6] = 7;
        layer_1_weights[90][6] = 6;
        layer_1_weights[91][6] = 5;
        layer_1_weights[92][6] = 0;
        layer_1_weights[93][6] = 3;
        layer_1_weights[94][6] = -4;
        layer_1_weights[95][6] = -6;
        layer_1_weights[96][6] = -14;
        layer_1_weights[97][6] = -7;
        layer_1_weights[98][6] = -17;
        layer_1_weights[99][6] = -15;
        layer_1_weights[100][6] = -18;
        layer_1_weights[101][6] = -9;
        layer_1_weights[102][6] = -3;
        layer_1_weights[103][6] = 1;
        layer_1_weights[104][6] = -2;
        layer_1_weights[105][6] = -5;
        layer_1_weights[106][6] = 1;
        layer_1_weights[107][6] = 9;
        layer_1_weights[108][6] = -7;
        layer_1_weights[109][6] = -3;
        layer_1_weights[110][6] = -13;
        layer_1_weights[111][6] = -8;
        layer_1_weights[112][6] = -10;
        layer_1_weights[113][6] = -4;
        layer_1_weights[114][6] = -4;
        layer_1_weights[115][6] = -2;
        layer_1_weights[116][6] = -5;
        layer_1_weights[117][6] = 0;
        layer_1_weights[118][6] = 5;
        layer_1_weights[119][6] = 11;
        layer_1_weights[120][6] = 2;
        layer_1_weights[121][6] = 14;
        layer_1_weights[122][6] = 14;
        layer_1_weights[123][6] = 6;
        layer_1_weights[124][6] = 5;
        layer_1_weights[125][6] = -2;
        layer_1_weights[126][6] = 0;
        layer_1_weights[127][6] = -4;
        layer_1_weights[128][6] = -5;
        layer_1_weights[129][6] = 2;
        layer_1_weights[130][6] = 11;
        layer_1_weights[131][6] = -3;
        layer_1_weights[132][6] = 0;
        layer_1_weights[133][6] = 9;
        layer_1_weights[134][6] = 4;
        layer_1_weights[135][6] = 11;
        layer_1_weights[136][6] = 9;
        layer_1_weights[137][6] = 9;
        layer_1_weights[138][6] = 18;
        layer_1_weights[139][6] = 10;
        layer_1_weights[140][6] = 12;
        layer_1_weights[141][6] = 11;
        layer_1_weights[142][6] = -2;
        layer_1_weights[143][6] = -1;
        layer_1_weights[0][7] = -3;
        layer_1_weights[1][7] = -1;
        layer_1_weights[2][7] = 1;
        layer_1_weights[3][7] = -4;
        layer_1_weights[4][7] = 4;
        layer_1_weights[5][7] = 11;
        layer_1_weights[6][7] = 9;
        layer_1_weights[7][7] = -10;
        layer_1_weights[8][7] = 1;
        layer_1_weights[9][7] = -12;
        layer_1_weights[10][7] = -1;
        layer_1_weights[11][7] = -2;
        layer_1_weights[12][7] = 2;
        layer_1_weights[13][7] = 3;
        layer_1_weights[14][7] = -7;
        layer_1_weights[15][7] = 0;
        layer_1_weights[16][7] = -12;
        layer_1_weights[17][7] = -5;
        layer_1_weights[18][7] = -5;
        layer_1_weights[19][7] = -4;
        layer_1_weights[20][7] = -1;
        layer_1_weights[21][7] = 1;
        layer_1_weights[22][7] = -7;
        layer_1_weights[23][7] = 3;
        layer_1_weights[24][7] = 1;
        layer_1_weights[25][7] = -3;
        layer_1_weights[26][7] = -3;
        layer_1_weights[27][7] = -8;
        layer_1_weights[28][7] = 0;
        layer_1_weights[29][7] = 4;
        layer_1_weights[30][7] = 10;
        layer_1_weights[31][7] = 9;
        layer_1_weights[32][7] = 4;
        layer_1_weights[33][7] = 4;
        layer_1_weights[34][7] = -4;
        layer_1_weights[35][7] = -1;
        layer_1_weights[36][7] = -8;
        layer_1_weights[37][7] = 4;
        layer_1_weights[38][7] = -3;
        layer_1_weights[39][7] = -4;
        layer_1_weights[40][7] = 6;
        layer_1_weights[41][7] = 14;
        layer_1_weights[42][7] = 12;
        layer_1_weights[43][7] = 12;
        layer_1_weights[44][7] = 8;
        layer_1_weights[45][7] = 5;
        layer_1_weights[46][7] = 14;
        layer_1_weights[47][7] = -15;
        layer_1_weights[48][7] = -10;
        layer_1_weights[49][7] = -14;
        layer_1_weights[50][7] = -3;
        layer_1_weights[51][7] = 4;
        layer_1_weights[52][7] = 10;
        layer_1_weights[53][7] = 2;
        layer_1_weights[54][7] = -11;
        layer_1_weights[55][7] = -3;
        layer_1_weights[56][7] = 4;
        layer_1_weights[57][7] = 3;
        layer_1_weights[58][7] = 5;
        layer_1_weights[59][7] = -5;
        layer_1_weights[60][7] = -2;
        layer_1_weights[61][7] = -2;
        layer_1_weights[62][7] = 4;
        layer_1_weights[63][7] = 4;
        layer_1_weights[64][7] = 6;
        layer_1_weights[65][7] = -1;
        layer_1_weights[66][7] = -13;
        layer_1_weights[67][7] = -5;
        layer_1_weights[68][7] = 3;
        layer_1_weights[69][7] = 9;
        layer_1_weights[70][7] = 10;
        layer_1_weights[71][7] = -4;
        layer_1_weights[72][7] = -9;
        layer_1_weights[73][7] = -4;
        layer_1_weights[74][7] = 2;
        layer_1_weights[75][7] = 4;
        layer_1_weights[76][7] = -2;
        layer_1_weights[77][7] = 2;
        layer_1_weights[78][7] = -11;
        layer_1_weights[79][7] = -3;
        layer_1_weights[80][7] = 2;
        layer_1_weights[81][7] = 6;
        layer_1_weights[82][7] = 11;
        layer_1_weights[83][7] = -3;
        layer_1_weights[84][7] = -16;
        layer_1_weights[85][7] = -8;
        layer_1_weights[86][7] = 9;
        layer_1_weights[87][7] = 10;
        layer_1_weights[88][7] = -2;
        layer_1_weights[89][7] = -6;
        layer_1_weights[90][7] = -5;
        layer_1_weights[91][7] = 0;
        layer_1_weights[92][7] = -6;
        layer_1_weights[93][7] = -4;
        layer_1_weights[94][7] = 1;
        layer_1_weights[95][7] = -4;
        layer_1_weights[96][7] = 15;
        layer_1_weights[97][7] = -5;
        layer_1_weights[98][7] = -1;
        layer_1_weights[99][7] = 7;
        layer_1_weights[100][7] = -1;
        layer_1_weights[101][7] = -3;
        layer_1_weights[102][7] = 0;
        layer_1_weights[103][7] = -3;
        layer_1_weights[104][7] = -6;
        layer_1_weights[105][7] = -1;
        layer_1_weights[106][7] = 1;
        layer_1_weights[107][7] = -4;
        layer_1_weights[108][7] = -12;
        layer_1_weights[109][7] = 0;
        layer_1_weights[110][7] = 5;
        layer_1_weights[111][7] = 3;
        layer_1_weights[112][7] = 8;
        layer_1_weights[113][7] = 3;
        layer_1_weights[114][7] = -6;
        layer_1_weights[115][7] = -8;
        layer_1_weights[116][7] = -4;
        layer_1_weights[117][7] = -1;
        layer_1_weights[118][7] = 6;
        layer_1_weights[119][7] = 0;
        layer_1_weights[120][7] = 1;
        layer_1_weights[121][7] = -7;
        layer_1_weights[122][7] = -2;
        layer_1_weights[123][7] = 3;
        layer_1_weights[124][7] = 4;
        layer_1_weights[125][7] = 3;
        layer_1_weights[126][7] = 5;
        layer_1_weights[127][7] = 5;
        layer_1_weights[128][7] = -2;
        layer_1_weights[129][7] = 6;
        layer_1_weights[130][7] = -2;
        layer_1_weights[131][7] = -9;
        layer_1_weights[132][7] = -1;
        layer_1_weights[133][7] = 4;
        layer_1_weights[134][7] = -4;
        layer_1_weights[135][7] = -3;
        layer_1_weights[136][7] = -4;
        layer_1_weights[137][7] = -3;
        layer_1_weights[138][7] = -1;
        layer_1_weights[139][7] = -2;
        layer_1_weights[140][7] = -6;
        layer_1_weights[141][7] = -9;
        layer_1_weights[142][7] = 1;
        layer_1_weights[143][7] = 2;
        layer_1_weights[0][8] = -1;
        layer_1_weights[1][8] = -2;
        layer_1_weights[2][8] = 0;
        layer_1_weights[3][8] = -5;
        layer_1_weights[4][8] = 2;
        layer_1_weights[5][8] = 2;
        layer_1_weights[6][8] = -6;
        layer_1_weights[7][8] = 1;
        layer_1_weights[8][8] = -1;
        layer_1_weights[9][8] = -6;
        layer_1_weights[10][8] = 0;
        layer_1_weights[11][8] = 2;
        layer_1_weights[12][8] = -3;
        layer_1_weights[13][8] = 1;
        layer_1_weights[14][8] = 1;
        layer_1_weights[15][8] = 1;
        layer_1_weights[16][8] = 2;
        layer_1_weights[17][8] = 2;
        layer_1_weights[18][8] = -4;
        layer_1_weights[19][8] = 0;
        layer_1_weights[20][8] = 1;
        layer_1_weights[21][8] = -3;
        layer_1_weights[22][8] = 11;
        layer_1_weights[23][8] = 10;
        layer_1_weights[24][8] = 1;
        layer_1_weights[25][8] = 11;
        layer_1_weights[26][8] = 8;
        layer_1_weights[27][8] = 14;
        layer_1_weights[28][8] = 10;
        layer_1_weights[29][8] = 9;
        layer_1_weights[30][8] = 2;
        layer_1_weights[31][8] = 1;
        layer_1_weights[32][8] = -1;
        layer_1_weights[33][8] = 0;
        layer_1_weights[34][8] = -1;
        layer_1_weights[35][8] = 16;
        layer_1_weights[36][8] = 9;
        layer_1_weights[37][8] = 17;
        layer_1_weights[38][8] = 8;
        layer_1_weights[39][8] = 9;
        layer_1_weights[40][8] = 7;
        layer_1_weights[41][8] = 6;
        layer_1_weights[42][8] = 3;
        layer_1_weights[43][8] = 6;
        layer_1_weights[44][8] = 1;
        layer_1_weights[45][8] = -2;
        layer_1_weights[46][8] = 2;
        layer_1_weights[47][8] = 7;
        layer_1_weights[48][8] = 2;
        layer_1_weights[49][8] = 16;
        layer_1_weights[50][8] = 5;
        layer_1_weights[51][8] = 4;
        layer_1_weights[52][8] = 3;
        layer_1_weights[53][8] = 5;
        layer_1_weights[54][8] = 1;
        layer_1_weights[55][8] = 4;
        layer_1_weights[56][8] = 2;
        layer_1_weights[57][8] = 1;
        layer_1_weights[58][8] = 10;
        layer_1_weights[59][8] = 0;
        layer_1_weights[60][8] = 24;
        layer_1_weights[61][8] = -5;
        layer_1_weights[62][8] = -9;
        layer_1_weights[63][8] = -11;
        layer_1_weights[64][8] = -6;
        layer_1_weights[65][8] = -5;
        layer_1_weights[66][8] = -11;
        layer_1_weights[67][8] = -1;
        layer_1_weights[68][8] = 3;
        layer_1_weights[69][8] = 0;
        layer_1_weights[70][8] = -2;
        layer_1_weights[71][8] = -17;
        layer_1_weights[72][8] = -1;
        layer_1_weights[73][8] = -34;
        layer_1_weights[74][8] = -23;
        layer_1_weights[75][8] = -9;
        layer_1_weights[76][8] = -6;
        layer_1_weights[77][8] = -3;
        layer_1_weights[78][8] = -2;
        layer_1_weights[79][8] = -1;
        layer_1_weights[80][8] = -1;
        layer_1_weights[81][8] = -6;
        layer_1_weights[82][8] = -4;
        layer_1_weights[83][8] = 3;
        layer_1_weights[84][8] = -3;
        layer_1_weights[85][8] = -25;
        layer_1_weights[86][8] = -4;
        layer_1_weights[87][8] = -1;
        layer_1_weights[88][8] = 4;
        layer_1_weights[89][8] = 4;
        layer_1_weights[90][8] = -5;
        layer_1_weights[91][8] = -1;
        layer_1_weights[92][8] = -2;
        layer_1_weights[93][8] = -1;
        layer_1_weights[94][8] = 0;
        layer_1_weights[95][8] = -3;
        layer_1_weights[96][8] = 20;
        layer_1_weights[97][8] = 7;
        layer_1_weights[98][8] = 6;
        layer_1_weights[99][8] = 0;
        layer_1_weights[100][8] = 2;
        layer_1_weights[101][8] = 0;
        layer_1_weights[102][8] = 1;
        layer_1_weights[103][8] = 1;
        layer_1_weights[104][8] = -2;
        layer_1_weights[105][8] = 2;
        layer_1_weights[106][8] = 1;
        layer_1_weights[107][8] = 0;
        layer_1_weights[108][8] = 13;
        layer_1_weights[109][8] = -3;
        layer_1_weights[110][8] = 4;
        layer_1_weights[111][8] = 6;
        layer_1_weights[112][8] = 6;
        layer_1_weights[113][8] = 8;
        layer_1_weights[114][8] = 8;
        layer_1_weights[115][8] = 3;
        layer_1_weights[116][8] = 5;
        layer_1_weights[117][8] = 5;
        layer_1_weights[118][8] = 2;
        layer_1_weights[119][8] = -11;
        layer_1_weights[120][8] = -2;
        layer_1_weights[121][8] = 4;
        layer_1_weights[122][8] = 3;
        layer_1_weights[123][8] = 6;
        layer_1_weights[124][8] = 7;
        layer_1_weights[125][8] = 7;
        layer_1_weights[126][8] = 5;
        layer_1_weights[127][8] = 3;
        layer_1_weights[128][8] = 4;
        layer_1_weights[129][8] = -4;
        layer_1_weights[130][8] = 6;
        layer_1_weights[131][8] = 10;
        layer_1_weights[132][8] = 3;
        layer_1_weights[133][8] = 11;
        layer_1_weights[134][8] = -7;
        layer_1_weights[135][8] = 11;
        layer_1_weights[136][8] = 14;
        layer_1_weights[137][8] = 9;
        layer_1_weights[138][8] = 11;
        layer_1_weights[139][8] = 13;
        layer_1_weights[140][8] = 15;
        layer_1_weights[141][8] = -2;
        layer_1_weights[142][8] = -2;
        layer_1_weights[143][8] = 3;
        layer_1_weights[0][9] = -1;
        layer_1_weights[1][9] = 3;
        layer_1_weights[2][9] = 1;
        layer_1_weights[3][9] = -4;
        layer_1_weights[4][9] = -12;
        layer_1_weights[5][9] = -23;
        layer_1_weights[6][9] = -2;
        layer_1_weights[7][9] = -4;
        layer_1_weights[8][9] = 0;
        layer_1_weights[9][9] = -4;
        layer_1_weights[10][9] = 0;
        layer_1_weights[11][9] = 0;
        layer_1_weights[12][9] = -2;
        layer_1_weights[13][9] = 1;
        layer_1_weights[14][9] = 10;
        layer_1_weights[15][9] = 11;
        layer_1_weights[16][9] = 8;
        layer_1_weights[17][9] = 4;
        layer_1_weights[18][9] = 0;
        layer_1_weights[19][9] = 3;
        layer_1_weights[20][9] = 0;
        layer_1_weights[21][9] = -4;
        layer_1_weights[22][9] = -2;
        layer_1_weights[23][9] = -4;
        layer_1_weights[24][9] = -3;
        layer_1_weights[25][9] = 2;
        layer_1_weights[26][9] = 11;
        layer_1_weights[27][9] = 4;
        layer_1_weights[28][9] = 7;
        layer_1_weights[29][9] = 7;
        layer_1_weights[30][9] = 5;
        layer_1_weights[31][9] = 6;
        layer_1_weights[32][9] = 2;
        layer_1_weights[33][9] = 6;
        layer_1_weights[34][9] = 4;
        layer_1_weights[35][9] = 0;
        layer_1_weights[36][9] = -3;
        layer_1_weights[37][9] = 12;
        layer_1_weights[38][9] = 5;
        layer_1_weights[39][9] = 4;
        layer_1_weights[40][9] = 5;
        layer_1_weights[41][9] = 0;
        layer_1_weights[42][9] = -1;
        layer_1_weights[43][9] = 1;
        layer_1_weights[44][9] = 0;
        layer_1_weights[45][9] = 1;
        layer_1_weights[46][9] = 2;
        layer_1_weights[47][9] = 9;
        layer_1_weights[48][9] = -7;
        layer_1_weights[49][9] = 6;
        layer_1_weights[50][9] = 0;
        layer_1_weights[51][9] = 3;
        layer_1_weights[52][9] = 4;
        layer_1_weights[53][9] = 1;
        layer_1_weights[54][9] = 1;
        layer_1_weights[55][9] = -1;
        layer_1_weights[56][9] = -3;
        layer_1_weights[57][9] = -6;
        layer_1_weights[58][9] = -5;
        layer_1_weights[59][9] = 5;
        layer_1_weights[60][9] = -24;
        layer_1_weights[61][9] = -8;
        layer_1_weights[62][9] = -9;
        layer_1_weights[63][9] = -5;
        layer_1_weights[64][9] = 4;
        layer_1_weights[65][9] = 18;
        layer_1_weights[66][9] = 15;
        layer_1_weights[67][9] = 7;
        layer_1_weights[68][9] = -1;
        layer_1_weights[69][9] = -2;
        layer_1_weights[70][9] = -8;
        layer_1_weights[71][9] = -4;
        layer_1_weights[72][9] = 12;
        layer_1_weights[73][9] = -19;
        layer_1_weights[74][9] = -18;
        layer_1_weights[75][9] = -15;
        layer_1_weights[76][9] = -8;
        layer_1_weights[77][9] = 8;
        layer_1_weights[78][9] = 6;
        layer_1_weights[79][9] = -1;
        layer_1_weights[80][9] = 2;
        layer_1_weights[81][9] = 2;
        layer_1_weights[82][9] = 7;
        layer_1_weights[83][9] = 13;
        layer_1_weights[84][9] = 16;
        layer_1_weights[85][9] = -2;
        layer_1_weights[86][9] = 0;
        layer_1_weights[87][9] = -11;
        layer_1_weights[88][9] = -29;
        layer_1_weights[89][9] = -18;
        layer_1_weights[90][9] = -1;
        layer_1_weights[91][9] = 2;
        layer_1_weights[92][9] = 3;
        layer_1_weights[93][9] = 1;
        layer_1_weights[94][9] = 6;
        layer_1_weights[95][9] = 10;
        layer_1_weights[96][9] = 16;
        layer_1_weights[97][9] = 9;
        layer_1_weights[98][9] = 10;
        layer_1_weights[99][9] = 7;
        layer_1_weights[100][9] = -6;
        layer_1_weights[101][9] = -1;
        layer_1_weights[102][9] = -1;
        layer_1_weights[103][9] = 2;
        layer_1_weights[104][9] = -1;
        layer_1_weights[105][9] = 4;
        layer_1_weights[106][9] = -3;
        layer_1_weights[107][9] = -2;
        layer_1_weights[108][9] = 6;
        layer_1_weights[109][9] = -1;
        layer_1_weights[110][9] = 0;
        layer_1_weights[111][9] = 5;
        layer_1_weights[112][9] = 4;
        layer_1_weights[113][9] = 1;
        layer_1_weights[114][9] = 1;
        layer_1_weights[115][9] = -1;
        layer_1_weights[116][9] = -1;
        layer_1_weights[117][9] = -4;
        layer_1_weights[118][9] = -9;
        layer_1_weights[119][9] = -10;
        layer_1_weights[120][9] = -1;
        layer_1_weights[121][9] = -2;
        layer_1_weights[122][9] = -2;
        layer_1_weights[123][9] = -1;
        layer_1_weights[124][9] = -4;
        layer_1_weights[125][9] = 0;
        layer_1_weights[126][9] = -1;
        layer_1_weights[127][9] = -3;
        layer_1_weights[128][9] = -2;
        layer_1_weights[129][9] = -11;
        layer_1_weights[130][9] = -15;
        layer_1_weights[131][9] = -4;
        layer_1_weights[132][9] = 1;
        layer_1_weights[133][9] = 11;
        layer_1_weights[134][9] = 0;
        layer_1_weights[135][9] = 8;
        layer_1_weights[136][9] = 6;
        layer_1_weights[137][9] = -1;
        layer_1_weights[138][9] = 7;
        layer_1_weights[139][9] = 3;
        layer_1_weights[140][9] = -9;
        layer_1_weights[141][9] = 5;
        layer_1_weights[142][9] = -1;
        layer_1_weights[143][9] = 1;
        layer_1_weights[0][10] = -3;
        layer_1_weights[1][10] = -2;
        layer_1_weights[2][10] = 4;
        layer_1_weights[3][10] = 11;
        layer_1_weights[4][10] = 18;
        layer_1_weights[5][10] = 5;
        layer_1_weights[6][10] = 3;
        layer_1_weights[7][10] = 8;
        layer_1_weights[8][10] = 8;
        layer_1_weights[9][10] = 4;
        layer_1_weights[10][10] = 3;
        layer_1_weights[11][10] = -2;
        layer_1_weights[12][10] = -1;
        layer_1_weights[13][10] = 2;
        layer_1_weights[14][10] = 8;
        layer_1_weights[15][10] = -2;
        layer_1_weights[16][10] = 0;
        layer_1_weights[17][10] = 1;
        layer_1_weights[18][10] = 1;
        layer_1_weights[19][10] = 1;
        layer_1_weights[20][10] = 3;
        layer_1_weights[21][10] = 2;
        layer_1_weights[22][10] = -1;
        layer_1_weights[23][10] = 6;
        layer_1_weights[24][10] = 2;
        layer_1_weights[25][10] = 11;
        layer_1_weights[26][10] = 1;
        layer_1_weights[27][10] = 0;
        layer_1_weights[28][10] = 1;
        layer_1_weights[29][10] = 8;
        layer_1_weights[30][10] = 16;
        layer_1_weights[31][10] = 7;
        layer_1_weights[32][10] = 5;
        layer_1_weights[33][10] = 4;
        layer_1_weights[34][10] = 4;
        layer_1_weights[35][10] = -1;
        layer_1_weights[36][10] = 8;
        layer_1_weights[37][10] = -6;
        layer_1_weights[38][10] = -8;
        layer_1_weights[39][10] = -3;
        layer_1_weights[40][10] = 8;
        layer_1_weights[41][10] = 10;
        layer_1_weights[42][10] = 7;
        layer_1_weights[43][10] = 9;
        layer_1_weights[44][10] = 4;
        layer_1_weights[45][10] = 3;
        layer_1_weights[46][10] = 0;
        layer_1_weights[47][10] = -5;
        layer_1_weights[48][10] = -1;
        layer_1_weights[49][10] = -8;
        layer_1_weights[50][10] = -10;
        layer_1_weights[51][10] = -8;
        layer_1_weights[52][10] = -8;
        layer_1_weights[53][10] = -23;
        layer_1_weights[54][10] = -12;
        layer_1_weights[55][10] = -4;
        layer_1_weights[56][10] = -1;
        layer_1_weights[57][10] = 4;
        layer_1_weights[58][10] = 2;
        layer_1_weights[59][10] = 0;
        layer_1_weights[60][10] = -10;
        layer_1_weights[61][10] = -6;
        layer_1_weights[62][10] = -5;
        layer_1_weights[63][10] = -3;
        layer_1_weights[64][10] = -9;
        layer_1_weights[65][10] = -8;
        layer_1_weights[66][10] = 3;
        layer_1_weights[67][10] = 7;
        layer_1_weights[68][10] = 0;
        layer_1_weights[69][10] = -3;
        layer_1_weights[70][10] = 4;
        layer_1_weights[71][10] = 8;
        layer_1_weights[72][10] = -11;
        layer_1_weights[73][10] = 2;
        layer_1_weights[74][10] = 9;
        layer_1_weights[75][10] = -3;
        layer_1_weights[76][10] = -2;
        layer_1_weights[77][10] = 3;
        layer_1_weights[78][10] = 10;
        layer_1_weights[79][10] = 0;
        layer_1_weights[80][10] = -3;
        layer_1_weights[81][10] = -6;
        layer_1_weights[82][10] = -10;
        layer_1_weights[83][10] = 6;
        layer_1_weights[84][10] = 2;
        layer_1_weights[85][10] = 5;
        layer_1_weights[86][10] = 2;
        layer_1_weights[87][10] = -1;
        layer_1_weights[88][10] = -3;
        layer_1_weights[89][10] = 1;
        layer_1_weights[90][10] = 3;
        layer_1_weights[91][10] = -3;
        layer_1_weights[92][10] = -4;
        layer_1_weights[93][10] = -14;
        layer_1_weights[94][10] = -18;
        layer_1_weights[95][10] = 1;
        layer_1_weights[96][10] = 2;
        layer_1_weights[97][10] = 0;
        layer_1_weights[98][10] = 8;
        layer_1_weights[99][10] = 7;
        layer_1_weights[100][10] = 3;
        layer_1_weights[101][10] = 8;
        layer_1_weights[102][10] = 3;
        layer_1_weights[103][10] = 0;
        layer_1_weights[104][10] = -1;
        layer_1_weights[105][10] = -4;
        layer_1_weights[106][10] = 9;
        layer_1_weights[107][10] = 13;
        layer_1_weights[108][10] = 12;
        layer_1_weights[109][10] = 6;
        layer_1_weights[110][10] = 2;
        layer_1_weights[111][10] = 3;
        layer_1_weights[112][10] = 2;
        layer_1_weights[113][10] = -3;
        layer_1_weights[114][10] = 1;
        layer_1_weights[115][10] = -5;
        layer_1_weights[116][10] = 5;
        layer_1_weights[117][10] = -1;
        layer_1_weights[118][10] = 5;
        layer_1_weights[119][10] = -9;
        layer_1_weights[120][10] = 1;
        layer_1_weights[121][10] = 1;
        layer_1_weights[122][10] = -4;
        layer_1_weights[123][10] = -10;
        layer_1_weights[124][10] = -9;
        layer_1_weights[125][10] = -6;
        layer_1_weights[126][10] = -3;
        layer_1_weights[127][10] = 1;
        layer_1_weights[128][10] = 5;
        layer_1_weights[129][10] = 4;
        layer_1_weights[130][10] = 16;
        layer_1_weights[131][10] = 14;
        layer_1_weights[132][10] = 1;
        layer_1_weights[133][10] = -1;
        layer_1_weights[134][10] = 1;
        layer_1_weights[135][10] = 3;
        layer_1_weights[136][10] = 5;
        layer_1_weights[137][10] = 1;
        layer_1_weights[138][10] = -1;
        layer_1_weights[139][10] = 10;
        layer_1_weights[140][10] = 5;
        layer_1_weights[141][10] = -2;
        layer_1_weights[142][10] = 3;
        layer_1_weights[143][10] = 0;
        layer_1_weights[0][11] = 1;
        layer_1_weights[1][11] = 3;
        layer_1_weights[2][11] = 7;
        layer_1_weights[3][11] = 17;
        layer_1_weights[4][11] = 22;
        layer_1_weights[5][11] = 13;
        layer_1_weights[6][11] = 18;
        layer_1_weights[7][11] = 9;
        layer_1_weights[8][11] = 10;
        layer_1_weights[9][11] = 16;
        layer_1_weights[10][11] = 1;
        layer_1_weights[11][11] = -3;
        layer_1_weights[12][11] = 2;
        layer_1_weights[13][11] = 2;
        layer_1_weights[14][11] = 10;
        layer_1_weights[15][11] = 2;
        layer_1_weights[16][11] = -8;
        layer_1_weights[17][11] = -6;
        layer_1_weights[18][11] = -7;
        layer_1_weights[19][11] = 0;
        layer_1_weights[20][11] = -4;
        layer_1_weights[21][11] = -11;
        layer_1_weights[22][11] = -17;
        layer_1_weights[23][11] = 12;
        layer_1_weights[24][11] = 1;
        layer_1_weights[25][11] = 5;
        layer_1_weights[26][11] = 2;
        layer_1_weights[27][11] = 6;
        layer_1_weights[28][11] = 2;
        layer_1_weights[29][11] = 1;
        layer_1_weights[30][11] = 0;
        layer_1_weights[31][11] = -5;
        layer_1_weights[32][11] = -1;
        layer_1_weights[33][11] = 0;
        layer_1_weights[34][11] = 4;
        layer_1_weights[35][11] = -7;
        layer_1_weights[36][11] = 19;
        layer_1_weights[37][11] = 5;
        layer_1_weights[38][11] = 0;
        layer_1_weights[39][11] = 4;
        layer_1_weights[40][11] = 0;
        layer_1_weights[41][11] = 3;
        layer_1_weights[42][11] = 1;
        layer_1_weights[43][11] = -4;
        layer_1_weights[44][11] = -3;
        layer_1_weights[45][11] = 4;
        layer_1_weights[46][11] = -4;
        layer_1_weights[47][11] = -2;
        layer_1_weights[48][11] = 6;
        layer_1_weights[49][11] = 9;
        layer_1_weights[50][11] = 5;
        layer_1_weights[51][11] = 1;
        layer_1_weights[52][11] = 0;
        layer_1_weights[53][11] = 1;
        layer_1_weights[54][11] = 1;
        layer_1_weights[55][11] = 1;
        layer_1_weights[56][11] = 0;
        layer_1_weights[57][11] = -1;
        layer_1_weights[58][11] = -8;
        layer_1_weights[59][11] = -1;
        layer_1_weights[60][11] = 13;
        layer_1_weights[61][11] = 7;
        layer_1_weights[62][11] = -1;
        layer_1_weights[63][11] = 7;
        layer_1_weights[64][11] = 2;
        layer_1_weights[65][11] = -6;
        layer_1_weights[66][11] = 2;
        layer_1_weights[67][11] = 5;
        layer_1_weights[68][11] = 3;
        layer_1_weights[69][11] = 1;
        layer_1_weights[70][11] = -3;
        layer_1_weights[71][11] = -4;
        layer_1_weights[72][11] = -3;
        layer_1_weights[73][11] = 3;
        layer_1_weights[74][11] = 5;
        layer_1_weights[75][11] = -4;
        layer_1_weights[76][11] = -10;
        layer_1_weights[77][11] = -11;
        layer_1_weights[78][11] = 10;
        layer_1_weights[79][11] = 2;
        layer_1_weights[80][11] = 1;
        layer_1_weights[81][11] = -5;
        layer_1_weights[82][11] = 5;
        layer_1_weights[83][11] = 10;
        layer_1_weights[84][11] = 1;
        layer_1_weights[85][11] = -15;
        layer_1_weights[86][11] = -4;
        layer_1_weights[87][11] = -14;
        layer_1_weights[88][11] = -17;
        layer_1_weights[89][11] = 6;
        layer_1_weights[90][11] = 10;
        layer_1_weights[91][11] = 5;
        layer_1_weights[92][11] = -1;
        layer_1_weights[93][11] = 0;
        layer_1_weights[94][11] = -6;
        layer_1_weights[95][11] = 7;
        layer_1_weights[96][11] = 2;
        layer_1_weights[97][11] = -25;
        layer_1_weights[98][11] = -8;
        layer_1_weights[99][11] = -21;
        layer_1_weights[100][11] = -5;
        layer_1_weights[101][11] = 18;
        layer_1_weights[102][11] = 9;
        layer_1_weights[103][11] = 4;
        layer_1_weights[104][11] = 3;
        layer_1_weights[105][11] = -3;
        layer_1_weights[106][11] = -5;
        layer_1_weights[107][11] = -4;
        layer_1_weights[108][11] = -2;
        layer_1_weights[109][11] = -1;
        layer_1_weights[110][11] = -12;
        layer_1_weights[111][11] = -1;
        layer_1_weights[112][11] = -8;
        layer_1_weights[113][11] = 4;
        layer_1_weights[114][11] = 5;
        layer_1_weights[115][11] = 3;
        layer_1_weights[116][11] = -1;
        layer_1_weights[117][11] = -4;
        layer_1_weights[118][11] = 0;
        layer_1_weights[119][11] = -1;
        layer_1_weights[120][11] = -3;
        layer_1_weights[121][11] = -13;
        layer_1_weights[122][11] = -13;
        layer_1_weights[123][11] = -11;
        layer_1_weights[124][11] = -11;
        layer_1_weights[125][11] = -7;
        layer_1_weights[126][11] = 0;
        layer_1_weights[127][11] = 2;
        layer_1_weights[128][11] = 2;
        layer_1_weights[129][11] = 5;
        layer_1_weights[130][11] = 3;
        layer_1_weights[131][11] = -2;
        layer_1_weights[132][11] = 1;
        layer_1_weights[133][11] = -1;
        layer_1_weights[134][11] = -18;
        layer_1_weights[135][11] = -1;
        layer_1_weights[136][11] = -1;
        layer_1_weights[137][11] = 1;
        layer_1_weights[138][11] = 4;
        layer_1_weights[139][11] = 5;
        layer_1_weights[140][11] = 3;
        layer_1_weights[141][11] = -5;
        layer_1_weights[142][11] = 2;
        layer_1_weights[143][11] = 1;
        layer_1_weights[0][12] = -3;
        layer_1_weights[1][12] = -1;
        layer_1_weights[2][12] = -8;
        layer_1_weights[3][12] = -12;
        layer_1_weights[4][12] = 6;
        layer_1_weights[5][12] = 1;
        layer_1_weights[6][12] = 5;
        layer_1_weights[7][12] = -2;
        layer_1_weights[8][12] = -3;
        layer_1_weights[9][12] = -18;
        layer_1_weights[10][12] = -1;
        layer_1_weights[11][12] = 2;
        layer_1_weights[12][12] = 2;
        layer_1_weights[13][12] = -1;
        layer_1_weights[14][12] = 2;
        layer_1_weights[15][12] = 0;
        layer_1_weights[16][12] = 6;
        layer_1_weights[17][12] = 3;
        layer_1_weights[18][12] = 11;
        layer_1_weights[19][12] = 13;
        layer_1_weights[20][12] = 0;
        layer_1_weights[21][12] = -2;
        layer_1_weights[22][12] = -12;
        layer_1_weights[23][12] = -6;
        layer_1_weights[24][12] = -2;
        layer_1_weights[25][12] = -8;
        layer_1_weights[26][12] = 7;
        layer_1_weights[27][12] = 1;
        layer_1_weights[28][12] = -2;
        layer_1_weights[29][12] = 4;
        layer_1_weights[30][12] = 3;
        layer_1_weights[31][12] = -3;
        layer_1_weights[32][12] = 4;
        layer_1_weights[33][12] = 4;
        layer_1_weights[34][12] = 4;
        layer_1_weights[35][12] = -11;
        layer_1_weights[36][12] = 4;
        layer_1_weights[37][12] = 15;
        layer_1_weights[38][12] = 4;
        layer_1_weights[39][12] = -2;
        layer_1_weights[40][12] = -6;
        layer_1_weights[41][12] = -9;
        layer_1_weights[42][12] = -5;
        layer_1_weights[43][12] = 6;
        layer_1_weights[44][12] = 11;
        layer_1_weights[45][12] = 8;
        layer_1_weights[46][12] = 17;
        layer_1_weights[47][12] = 5;
        layer_1_weights[48][12] = 8;
        layer_1_weights[49][12] = 2;
        layer_1_weights[50][12] = -10;
        layer_1_weights[51][12] = -10;
        layer_1_weights[52][12] = -8;
        layer_1_weights[53][12] = -8;
        layer_1_weights[54][12] = -3;
        layer_1_weights[55][12] = 9;
        layer_1_weights[56][12] = 9;
        layer_1_weights[57][12] = 9;
        layer_1_weights[58][12] = 5;
        layer_1_weights[59][12] = 3;
        layer_1_weights[60][12] = 5;
        layer_1_weights[61][12] = -12;
        layer_1_weights[62][12] = -4;
        layer_1_weights[63][12] = 5;
        layer_1_weights[64][12] = 7;
        layer_1_weights[65][12] = 4;
        layer_1_weights[66][12] = -9;
        layer_1_weights[67][12] = -2;
        layer_1_weights[68][12] = -4;
        layer_1_weights[69][12] = -7;
        layer_1_weights[70][12] = -16;
        layer_1_weights[71][12] = -5;
        layer_1_weights[72][12] = 11;
        layer_1_weights[73][12] = 9;
        layer_1_weights[74][12] = 13;
        layer_1_weights[75][12] = 10;
        layer_1_weights[76][12] = 5;
        layer_1_weights[77][12] = 3;
        layer_1_weights[78][12] = -5;
        layer_1_weights[79][12] = 2;
        layer_1_weights[80][12] = -3;
        layer_1_weights[81][12] = -3;
        layer_1_weights[82][12] = 4;
        layer_1_weights[83][12] = -16;
        layer_1_weights[84][12] = 17;
        layer_1_weights[85][12] = 11;
        layer_1_weights[86][12] = 9;
        layer_1_weights[87][12] = 1;
        layer_1_weights[88][12] = -3;
        layer_1_weights[89][12] = 0;
        layer_1_weights[90][12] = 6;
        layer_1_weights[91][12] = 4;
        layer_1_weights[92][12] = 0;
        layer_1_weights[93][12] = 2;
        layer_1_weights[94][12] = 0;
        layer_1_weights[95][12] = -2;
        layer_1_weights[96][12] = 24;
        layer_1_weights[97][12] = 7;
        layer_1_weights[98][12] = 7;
        layer_1_weights[99][12] = 2;
        layer_1_weights[100][12] = -4;
        layer_1_weights[101][12] = -2;
        layer_1_weights[102][12] = 1;
        layer_1_weights[103][12] = 4;
        layer_1_weights[104][12] = 3;
        layer_1_weights[105][12] = -4;
        layer_1_weights[106][12] = -6;
        layer_1_weights[107][12] = -3;
        layer_1_weights[108][12] = 13;
        layer_1_weights[109][12] = 4;
        layer_1_weights[110][12] = 0;
        layer_1_weights[111][12] = -1;
        layer_1_weights[112][12] = -3;
        layer_1_weights[113][12] = -3;
        layer_1_weights[114][12] = -3;
        layer_1_weights[115][12] = 3;
        layer_1_weights[116][12] = 9;
        layer_1_weights[117][12] = 3;
        layer_1_weights[118][12] = 11;
        layer_1_weights[119][12] = 2;
        layer_1_weights[120][12] = 2;
        layer_1_weights[121][12] = 5;
        layer_1_weights[122][12] = 5;
        layer_1_weights[123][12] = 5;
        layer_1_weights[124][12] = 3;
        layer_1_weights[125][12] = 4;
        layer_1_weights[126][12] = -2;
        layer_1_weights[127][12] = 0;
        layer_1_weights[128][12] = 0;
        layer_1_weights[129][12] = 1;
        layer_1_weights[130][12] = -1;
        layer_1_weights[131][12] = 3;
        layer_1_weights[132][12] = -2;
        layer_1_weights[133][12] = -1;
        layer_1_weights[134][12] = -3;
        layer_1_weights[135][12] = -2;
        layer_1_weights[136][12] = -3;
        layer_1_weights[137][12] = 0;
        layer_1_weights[138][12] = 0;
        layer_1_weights[139][12] = -1;
        layer_1_weights[140][12] = -6;
        layer_1_weights[141][12] = -10;
        layer_1_weights[142][12] = -1;
        layer_1_weights[143][12] = -1;
        layer_1_weights[0][13] = 2;
        layer_1_weights[1][13] = 2;
        layer_1_weights[2][13] = 4;
        layer_1_weights[3][13] = 20;
        layer_1_weights[4][13] = 16;
        layer_1_weights[5][13] = 15;
        layer_1_weights[6][13] = 2;
        layer_1_weights[7][13] = 23;
        layer_1_weights[8][13] = 3;
        layer_1_weights[9][13] = 22;
        layer_1_weights[10][13] = 1;
        layer_1_weights[11][13] = 0;
        layer_1_weights[12][13] = -2;
        layer_1_weights[13][13] = -2;
        layer_1_weights[14][13] = -2;
        layer_1_weights[15][13] = 1;
        layer_1_weights[16][13] = 2;
        layer_1_weights[17][13] = -8;
        layer_1_weights[18][13] = -4;
        layer_1_weights[19][13] = 5;
        layer_1_weights[20][13] = 9;
        layer_1_weights[21][13] = 6;
        layer_1_weights[22][13] = -2;
        layer_1_weights[23][13] = 5;
        layer_1_weights[24][13] = 1;
        layer_1_weights[25][13] = 8;
        layer_1_weights[26][13] = 9;
        layer_1_weights[27][13] = 2;
        layer_1_weights[28][13] = -3;
        layer_1_weights[29][13] = -3;
        layer_1_weights[30][13] = -3;
        layer_1_weights[31][13] = 1;
        layer_1_weights[32][13] = 4;
        layer_1_weights[33][13] = 5;
        layer_1_weights[34][13] = 11;
        layer_1_weights[35][13] = 11;
        layer_1_weights[36][13] = 16;
        layer_1_weights[37][13] = 12;
        layer_1_weights[38][13] = 5;
        layer_1_weights[39][13] = 9;
        layer_1_weights[40][13] = 3;
        layer_1_weights[41][13] = -10;
        layer_1_weights[42][13] = -5;
        layer_1_weights[43][13] = 0;
        layer_1_weights[44][13] = 1;
        layer_1_weights[45][13] = 2;
        layer_1_weights[46][13] = 2;
        layer_1_weights[47][13] = 3;
        layer_1_weights[48][13] = 16;
        layer_1_weights[49][13] = 20;
        layer_1_weights[50][13] = 4;
        layer_1_weights[51][13] = 5;
        layer_1_weights[52][13] = 0;
        layer_1_weights[53][13] = 1;
        layer_1_weights[54][13] = 1;
        layer_1_weights[55][13] = -2;
        layer_1_weights[56][13] = 0;
        layer_1_weights[57][13] = -1;
        layer_1_weights[58][13] = 0;
        layer_1_weights[59][13] = -4;
        layer_1_weights[60][13] = 9;
        layer_1_weights[61][13] = -8;
        layer_1_weights[62][13] = 4;
        layer_1_weights[63][13] = 6;
        layer_1_weights[64][13] = 5;
        layer_1_weights[65][13] = 6;
        layer_1_weights[66][13] = 6;
        layer_1_weights[67][13] = 3;
        layer_1_weights[68][13] = 2;
        layer_1_weights[69][13] = 5;
        layer_1_weights[70][13] = 4;
        layer_1_weights[71][13] = -9;
        layer_1_weights[72][13] = -1;
        layer_1_weights[73][13] = 0;
        layer_1_weights[74][13] = 3;
        layer_1_weights[75][13] = -3;
        layer_1_weights[76][13] = 3;
        layer_1_weights[77][13] = -4;
        layer_1_weights[78][13] = -8;
        layer_1_weights[79][13] = -5;
        layer_1_weights[80][13] = 8;
        layer_1_weights[81][13] = 8;
        layer_1_weights[82][13] = 8;
        layer_1_weights[83][13] = -13;
        layer_1_weights[84][13] = 13;
        layer_1_weights[85][13] = 0;
        layer_1_weights[86][13] = 0;
        layer_1_weights[87][13] = 4;
        layer_1_weights[88][13] = -4;
        layer_1_weights[89][13] = -4;
        layer_1_weights[90][13] = -9;
        layer_1_weights[91][13] = 5;
        layer_1_weights[92][13] = 6;
        layer_1_weights[93][13] = -3;
        layer_1_weights[94][13] = 3;
        layer_1_weights[95][13] = -8;
        layer_1_weights[96][13] = 14;
        layer_1_weights[97][13] = 10;
        layer_1_weights[98][13] = -7;
        layer_1_weights[99][13] = -5;
        layer_1_weights[100][13] = 4;
        layer_1_weights[101][13] = 4;
        layer_1_weights[102][13] = 1;
        layer_1_weights[103][13] = 12;
        layer_1_weights[104][13] = 2;
        layer_1_weights[105][13] = -3;
        layer_1_weights[106][13] = -9;
        layer_1_weights[107][13] = -26;
        layer_1_weights[108][13] = 7;
        layer_1_weights[109][13] = -15;
        layer_1_weights[110][13] = -11;
        layer_1_weights[111][13] = -4;
        layer_1_weights[112][13] = 3;
        layer_1_weights[113][13] = 10;
        layer_1_weights[114][13] = 8;
        layer_1_weights[115][13] = 3;
        layer_1_weights[116][13] = -4;
        layer_1_weights[117][13] = -11;
        layer_1_weights[118][13] = -9;
        layer_1_weights[119][13] = 12;
        layer_1_weights[120][13] = 2;
        layer_1_weights[121][13] = 3;
        layer_1_weights[122][13] = -3;
        layer_1_weights[123][13] = -8;
        layer_1_weights[124][13] = -6;
        layer_1_weights[125][13] = 6;
        layer_1_weights[126][13] = 7;
        layer_1_weights[127][13] = -1;
        layer_1_weights[128][13] = -6;
        layer_1_weights[129][13] = -7;
        layer_1_weights[130][13] = -13;
        layer_1_weights[131][13] = -2;
        layer_1_weights[132][13] = 2;
        layer_1_weights[133][13] = 1;
        layer_1_weights[134][13] = -2;
        layer_1_weights[135][13] = 9;
        layer_1_weights[136][13] = 9;
        layer_1_weights[137][13] = 3;
        layer_1_weights[138][13] = -2;
        layer_1_weights[139][13] = -5;
        layer_1_weights[140][13] = 5;
        layer_1_weights[141][13] = 10;
        layer_1_weights[142][13] = 2;
        layer_1_weights[143][13] = -2;
        layer_1_weights[0][14] = 0;
        layer_1_weights[1][14] = 1;
        layer_1_weights[2][14] = 2;
        layer_1_weights[3][14] = 11;
        layer_1_weights[4][14] = 4;
        layer_1_weights[5][14] = 0;
        layer_1_weights[6][14] = 11;
        layer_1_weights[7][14] = 0;
        layer_1_weights[8][14] = -17;
        layer_1_weights[9][14] = -3;
        layer_1_weights[10][14] = -1;
        layer_1_weights[11][14] = 0;
        layer_1_weights[12][14] = 1;
        layer_1_weights[13][14] = 0;
        layer_1_weights[14][14] = 8;
        layer_1_weights[15][14] = 1;
        layer_1_weights[16][14] = 0;
        layer_1_weights[17][14] = 3;
        layer_1_weights[18][14] = 4;
        layer_1_weights[19][14] = 1;
        layer_1_weights[20][14] = -1;
        layer_1_weights[21][14] = -11;
        layer_1_weights[22][14] = -16;
        layer_1_weights[23][14] = 11;
        layer_1_weights[24][14] = 3;
        layer_1_weights[25][14] = 2;
        layer_1_weights[26][14] = -6;
        layer_1_weights[27][14] = -9;
        layer_1_weights[28][14] = -9;
        layer_1_weights[29][14] = -9;
        layer_1_weights[30][14] = -6;
        layer_1_weights[31][14] = 9;
        layer_1_weights[32][14] = -4;
        layer_1_weights[33][14] = 3;
        layer_1_weights[34][14] = -3;
        layer_1_weights[35][14] = 1;
        layer_1_weights[36][14] = 8;
        layer_1_weights[37][14] = 1;
        layer_1_weights[38][14] = -1;
        layer_1_weights[39][14] = 1;
        layer_1_weights[40][14] = -1;
        layer_1_weights[41][14] = -9;
        layer_1_weights[42][14] = 4;
        layer_1_weights[43][14] = 9;
        layer_1_weights[44][14] = 1;
        layer_1_weights[45][14] = 0;
        layer_1_weights[46][14] = -3;
        layer_1_weights[47][14] = -11;
        layer_1_weights[48][14] = -3;
        layer_1_weights[49][14] = -2;
        layer_1_weights[50][14] = 8;
        layer_1_weights[51][14] = 9;
        layer_1_weights[52][14] = 3;
        layer_1_weights[53][14] = -6;
        layer_1_weights[54][14] = 8;
        layer_1_weights[55][14] = 4;
        layer_1_weights[56][14] = -3;
        layer_1_weights[57][14] = -3;
        layer_1_weights[58][14] = -11;
        layer_1_weights[59][14] = 4;
        layer_1_weights[60][14] = 6;
        layer_1_weights[61][14] = 8;
        layer_1_weights[62][14] = 6;
        layer_1_weights[63][14] = 7;
        layer_1_weights[64][14] = -9;
        layer_1_weights[65][14] = -7;
        layer_1_weights[66][14] = 11;
        layer_1_weights[67][14] = 1;
        layer_1_weights[68][14] = -4;
        layer_1_weights[69][14] = 2;
        layer_1_weights[70][14] = 3;
        layer_1_weights[71][14] = -1;
        layer_1_weights[72][14] = 4;
        layer_1_weights[73][14] = 5;
        layer_1_weights[74][14] = -8;
        layer_1_weights[75][14] = -15;
        layer_1_weights[76][14] = -5;
        layer_1_weights[77][14] = 13;
        layer_1_weights[78][14] = 6;
        layer_1_weights[79][14] = -5;
        layer_1_weights[80][14] = -3;
        layer_1_weights[81][14] = -8;
        layer_1_weights[82][14] = -11;
        layer_1_weights[83][14] = 5;
        layer_1_weights[84][14] = 0;
        layer_1_weights[85][14] = -2;
        layer_1_weights[86][14] = -18;
        layer_1_weights[87][14] = -2;
        layer_1_weights[88][14] = 6;
        layer_1_weights[89][14] = 7;
        layer_1_weights[90][14] = -5;
        layer_1_weights[91][14] = -9;
        layer_1_weights[92][14] = -7;
        layer_1_weights[93][14] = -13;
        layer_1_weights[94][14] = 2;
        layer_1_weights[95][14] = 18;
        layer_1_weights[96][14] = -4;
        layer_1_weights[97][14] = -5;
        layer_1_weights[98][14] = -4;
        layer_1_weights[99][14] = 5;
        layer_1_weights[100][14] = 9;
        layer_1_weights[101][14] = 3;
        layer_1_weights[102][14] = -5;
        layer_1_weights[103][14] = 4;
        layer_1_weights[104][14] = 6;
        layer_1_weights[105][14] = 10;
        layer_1_weights[106][14] = 11;
        layer_1_weights[107][14] = 33;
        layer_1_weights[108][14] = 2;
        layer_1_weights[109][14] = -5;
        layer_1_weights[110][14] = 3;
        layer_1_weights[111][14] = -2;
        layer_1_weights[112][14] = 3;
        layer_1_weights[113][14] = -1;
        layer_1_weights[114][14] = 2;
        layer_1_weights[115][14] = 5;
        layer_1_weights[116][14] = 8;
        layer_1_weights[117][14] = 5;
        layer_1_weights[118][14] = -3;
        layer_1_weights[119][14] = 5;
        layer_1_weights[120][14] = 2;
        layer_1_weights[121][14] = -9;
        layer_1_weights[122][14] = -1;
        layer_1_weights[123][14] = -4;
        layer_1_weights[124][14] = -2;
        layer_1_weights[125][14] = 0;
        layer_1_weights[126][14] = 0;
        layer_1_weights[127][14] = -7;
        layer_1_weights[128][14] = -4;
        layer_1_weights[129][14] = -4;
        layer_1_weights[130][14] = -1;
        layer_1_weights[131][14] = 15;
        layer_1_weights[132][14] = 2;
        layer_1_weights[133][14] = -15;
        layer_1_weights[134][14] = 9;
        layer_1_weights[135][14] = 1;
        layer_1_weights[136][14] = -1;
        layer_1_weights[137][14] = -12;
        layer_1_weights[138][14] = -7;
        layer_1_weights[139][14] = -20;
        layer_1_weights[140][14] = -14;
        layer_1_weights[141][14] = -8;
        layer_1_weights[142][14] = 0;
        layer_1_weights[143][14] = 3;
        layer_1_weights[0][15] = 3;
        layer_1_weights[1][15] = 2;
        layer_1_weights[2][15] = -1;
        layer_1_weights[3][15] = -10;
        layer_1_weights[4][15] = -18;
        layer_1_weights[5][15] = 0;
        layer_1_weights[6][15] = 6;
        layer_1_weights[7][15] = -4;
        layer_1_weights[8][15] = 13;
        layer_1_weights[9][15] = -19;
        layer_1_weights[10][15] = 2;
        layer_1_weights[11][15] = -3;
        layer_1_weights[12][15] = -1;
        layer_1_weights[13][15] = -3;
        layer_1_weights[14][15] = 22;
        layer_1_weights[15][15] = 0;
        layer_1_weights[16][15] = -4;
        layer_1_weights[17][15] = 0;
        layer_1_weights[18][15] = -9;
        layer_1_weights[19][15] = -11;
        layer_1_weights[20][15] = -7;
        layer_1_weights[21][15] = -5;
        layer_1_weights[22][15] = -2;
        layer_1_weights[23][15] = -7;
        layer_1_weights[24][15] = 0;
        layer_1_weights[25][15] = 20;
        layer_1_weights[26][15] = 11;
        layer_1_weights[27][15] = 11;
        layer_1_weights[28][15] = 7;
        layer_1_weights[29][15] = 3;
        layer_1_weights[30][15] = -3;
        layer_1_weights[31][15] = -5;
        layer_1_weights[32][15] = -7;
        layer_1_weights[33][15] = -8;
        layer_1_weights[34][15] = -10;
        layer_1_weights[35][15] = 1;
        layer_1_weights[36][15] = 14;
        layer_1_weights[37][15] = 17;
        layer_1_weights[38][15] = 11;
        layer_1_weights[39][15] = 5;
        layer_1_weights[40][15] = 1;
        layer_1_weights[41][15] = 3;
        layer_1_weights[42][15] = 9;
        layer_1_weights[43][15] = 5;
        layer_1_weights[44][15] = -6;
        layer_1_weights[45][15] = -3;
        layer_1_weights[46][15] = -11;
        layer_1_weights[47][15] = -5;
        layer_1_weights[48][15] = 13;
        layer_1_weights[49][15] = 3;
        layer_1_weights[50][15] = -4;
        layer_1_weights[51][15] = -7;
        layer_1_weights[52][15] = -6;
        layer_1_weights[53][15] = 0;
        layer_1_weights[54][15] = 7;
        layer_1_weights[55][15] = 7;
        layer_1_weights[56][15] = 2;
        layer_1_weights[57][15] = -8;
        layer_1_weights[58][15] = -13;
        layer_1_weights[59][15] = -6;
        layer_1_weights[60][15] = 27;
        layer_1_weights[61][15] = -4;
        layer_1_weights[62][15] = -9;
        layer_1_weights[63][15] = -7;
        layer_1_weights[64][15] = 3;
        layer_1_weights[65][15] = -3;
        layer_1_weights[66][15] = 6;
        layer_1_weights[67][15] = 10;
        layer_1_weights[68][15] = 3;
        layer_1_weights[69][15] = -4;
        layer_1_weights[70][15] = -19;
        layer_1_weights[71][15] = -18;
        layer_1_weights[72][15] = 20;
        layer_1_weights[73][15] = 8;
        layer_1_weights[74][15] = -4;
        layer_1_weights[75][15] = 1;
        layer_1_weights[76][15] = 5;
        layer_1_weights[77][15] = -3;
        layer_1_weights[78][15] = 12;
        layer_1_weights[79][15] = 11;
        layer_1_weights[80][15] = 4;
        layer_1_weights[81][15] = 1;
        layer_1_weights[82][15] = -7;
        layer_1_weights[83][15] = -10;
        layer_1_weights[84][15] = 11;
        layer_1_weights[85][15] = -4;
        layer_1_weights[86][15] = -6;
        layer_1_weights[87][15] = -4;
        layer_1_weights[88][15] = -2;
        layer_1_weights[89][15] = 1;
        layer_1_weights[90][15] = 6;
        layer_1_weights[91][15] = 2;
        layer_1_weights[92][15] = -2;
        layer_1_weights[93][15] = -2;
        layer_1_weights[94][15] = 1;
        layer_1_weights[95][15] = -3;
        layer_1_weights[96][15] = 10;
        layer_1_weights[97][15] = -5;
        layer_1_weights[98][15] = -3;
        layer_1_weights[99][15] = -6;
        layer_1_weights[100][15] = -7;
        layer_1_weights[101][15] = 1;
        layer_1_weights[102][15] = 3;
        layer_1_weights[103][15] = -7;
        layer_1_weights[104][15] = -6;
        layer_1_weights[105][15] = -3;
        layer_1_weights[106][15] = -8;
        layer_1_weights[107][15] = 0;
        layer_1_weights[108][15] = 9;
        layer_1_weights[109][15] = -1;
        layer_1_weights[110][15] = -2;
        layer_1_weights[111][15] = -1;
        layer_1_weights[112][15] = -1;
        layer_1_weights[113][15] = -1;
        layer_1_weights[114][15] = -3;
        layer_1_weights[115][15] = -2;
        layer_1_weights[116][15] = -2;
        layer_1_weights[117][15] = -4;
        layer_1_weights[118][15] = -17;
        layer_1_weights[119][15] = 0;
        layer_1_weights[120][15] = 3;
        layer_1_weights[121][15] = 16;
        layer_1_weights[122][15] = 5;
        layer_1_weights[123][15] = 4;
        layer_1_weights[124][15] = 3;
        layer_1_weights[125][15] = 1;
        layer_1_weights[126][15] = 0;
        layer_1_weights[127][15] = -2;
        layer_1_weights[128][15] = 1;
        layer_1_weights[129][15] = -8;
        layer_1_weights[130][15] = -5;
        layer_1_weights[131][15] = -1;
        layer_1_weights[132][15] = 0;
        layer_1_weights[133][15] = 14;
        layer_1_weights[134][15] = 16;
        layer_1_weights[135][15] = 11;
        layer_1_weights[136][15] = 2;
        layer_1_weights[137][15] = -3;
        layer_1_weights[138][15] = -4;
        layer_1_weights[139][15] = -10;
        layer_1_weights[140][15] = -4;
        layer_1_weights[141][15] = -10;
        layer_1_weights[142][15] = 2;
        layer_1_weights[143][15] = 3;
        layer_1_biases[0] = 5;
        layer_1_biases[1] = -9;
        layer_1_biases[2] = -16;
        layer_1_biases[3] = 4;
        layer_1_biases[4] = 2;
        layer_1_biases[5] = 12;
        layer_1_biases[6] = 11;
        layer_1_biases[7] = -2;
        layer_1_biases[8] = -19;
        layer_1_biases[9] = -5;
        layer_1_biases[10] = -8;
        layer_1_biases[11] = -3;
        layer_1_biases[12] = 3;
        layer_1_biases[13] = 4;
        layer_1_biases[14] = 1;
        layer_1_biases[15] = 8;
        layer_2_weights[0][0] = -4;
        layer_2_weights[1][0] = 4;
        layer_2_weights[2][0] = -2;
        layer_2_weights[3][0] = 0;
        layer_2_weights[4][0] = -14;
        layer_2_weights[5][0] = -9;
        layer_2_weights[6][0] = -18;
        layer_2_weights[7][0] = 17;
        layer_2_weights[8][0] = 1;
        layer_2_weights[9][0] = -28;
        layer_2_weights[10][0] = -21;
        layer_2_weights[11][0] = -5;
        layer_2_weights[12][0] = 5;
        layer_2_weights[13][0] = 11;
        layer_2_weights[14][0] = -5;
        layer_2_weights[15][0] = 9;
        layer_2_weights[0][1] = -3;
        layer_2_weights[1][1] = -20;
        layer_2_weights[2][1] = 6;
        layer_2_weights[3][1] = 12;
        layer_2_weights[4][1] = 7;
        layer_2_weights[5][1] = -13;
        layer_2_weights[6][1] = -18;
        layer_2_weights[7][1] = -23;
        layer_2_weights[8][1] = -20;
        layer_2_weights[9][1] = -2;
        layer_2_weights[10][1] = 1;
        layer_2_weights[11][1] = 18;
        layer_2_weights[12][1] = 3;
        layer_2_weights[13][1] = -21;
        layer_2_weights[14][1] = 19;
        layer_2_weights[15][1] = 1;
        layer_2_weights[0][2] = 24;
        layer_2_weights[1][2] = 0;
        layer_2_weights[2][2] = -9;
        layer_2_weights[3][2] = 3;
        layer_2_weights[4][2] = -10;
        layer_2_weights[5][2] = -26;
        layer_2_weights[6][2] = -6;
        layer_2_weights[7][2] = -4;
        layer_2_weights[8][2] = 24;
        layer_2_weights[9][2] = -11;
        layer_2_weights[10][2] = 9;
        layer_2_weights[11][2] = 4;
        layer_2_weights[12][2] = 16;
        layer_2_weights[13][2] = -16;
        layer_2_weights[14][2] = 16;
        layer_2_weights[15][2] = -7;
        layer_2_weights[0][3] = -5;
        layer_2_weights[1][3] = -4;
        layer_2_weights[2][3] = 7;
        layer_2_weights[3][3] = 7;
        layer_2_weights[4][3] = -14;
        layer_2_weights[5][3] = -10;
        layer_2_weights[6][3] = 5;
        layer_2_weights[7][3] = -13;
        layer_2_weights[8][3] = 5;
        layer_2_weights[9][3] = 11;
        layer_2_weights[10][3] = 11;
        layer_2_weights[11][3] = -19;
        layer_2_weights[12][3] = 10;
        layer_2_weights[13][3] = 1;
        layer_2_weights[14][3] = -11;
        layer_2_weights[15][3] = 2;
        layer_2_weights[0][4] = -9;
        layer_2_weights[1][4] = 10;
        layer_2_weights[2][4] = -12;
        layer_2_weights[3][4] = -29;
        layer_2_weights[4][4] = 13;
        layer_2_weights[5][4] = -25;
        layer_2_weights[6][4] = 3;
        layer_2_weights[7][4] = -3;
        layer_2_weights[8][4] = -14;
        layer_2_weights[9][4] = 9;
        layer_2_weights[10][4] = -33;
        layer_2_weights[11][4] = -10;
        layer_2_weights[12][4] = 12;
        layer_2_weights[13][4] = -6;
        layer_2_weights[14][4] = 5;
        layer_2_weights[15][4] = 12;
        layer_2_weights[0][5] = -5;
        layer_2_weights[1][5] = 3;
        layer_2_weights[2][5] = -6;
        layer_2_weights[3][5] = 17;
        layer_2_weights[4][5] = -1;
        layer_2_weights[5][5] = 29;
        layer_2_weights[6][5] = 5;
        layer_2_weights[7][5] = -10;
        layer_2_weights[8][5] = 0;
        layer_2_weights[9][5] = 8;
        layer_2_weights[10][5] = 8;
        layer_2_weights[11][5] = -23;
        layer_2_weights[12][5] = -16;
        layer_2_weights[13][5] = 5;
        layer_2_weights[14][5] = -21;
        layer_2_weights[15][5] = -20;
        layer_2_weights[0][6] = 16;
        layer_2_weights[1][6] = 11;
        layer_2_weights[2][6] = -6;
        layer_2_weights[3][6] = 9;
        layer_2_weights[4][6] = 5;
        layer_2_weights[5][6] = -6;
        layer_2_weights[6][6] = -37;
        layer_2_weights[7][6] = 0;
        layer_2_weights[8][6] = -18;
        layer_2_weights[9][6] = -31;
        layer_2_weights[10][6] = -10;
        layer_2_weights[11][6] = 14;
        layer_2_weights[12][6] = -17;
        layer_2_weights[13][6] = 11;
        layer_2_weights[14][6] = 0;
        layer_2_weights[15][6] = -3;
        layer_2_weights[0][7] = -6;
        layer_2_weights[1][7] = -21;
        layer_2_weights[2][7] = -14;
        layer_2_weights[3][7] = -20;
        layer_2_weights[4][7] = -8;
        layer_2_weights[5][7] = -2;
        layer_2_weights[6][7] = 18;
        layer_2_weights[7][7] = -1;
        layer_2_weights[8][7] = 6;
        layer_2_weights[9][7] = -10;
        layer_2_weights[10][7] = 14;
        layer_2_weights[11][7] = -5;
        layer_2_weights[12][7] = 0;
        layer_2_weights[13][7] = 6;
        layer_2_weights[14][7] = 6;
        layer_2_weights[15][7] = 14;
        layer_2_weights[0][8] = -13;
        layer_2_weights[1][8] = 5;
        layer_2_weights[2][8] = 17;
        layer_2_weights[3][8] = -8;
        layer_2_weights[4][8] = 11;
        layer_2_weights[5][8] = -5;
        layer_2_weights[6][8] = -11;
        layer_2_weights[7][8] = 1;
        layer_2_weights[8][8] = 9;
        layer_2_weights[9][8] = 6;
        layer_2_weights[10][8] = -1;
        layer_2_weights[11][8] = 11;
        layer_2_weights[12][8] = -5;
        layer_2_weights[13][8] = -6;
        layer_2_weights[14][8] = -4;
        layer_2_weights[15][8] = -18;
        layer_2_weights[0][9] = -35;
        layer_2_weights[1][9] = 12;
        layer_2_weights[2][9] = 8;
        layer_2_weights[3][9] = -14;
        layer_2_weights[4][9] = -10;
        layer_2_weights[5][9] = -3;
        layer_2_weights[6][9] = 9;
        layer_2_weights[7][9] = 9;
        layer_2_weights[8][9] = -21;
        layer_2_weights[9][9] = 20;
        layer_2_weights[10][9] = -2;
        layer_2_weights[11][9] = -12;
        layer_2_weights[12][9] = -13;
        layer_2_weights[13][9] = -6;
        layer_2_weights[14][9] = -23;
        layer_2_weights[15][9] = 10;
        layer_2_biases[0] = -5;
        layer_2_biases[1] = 14;
        layer_2_biases[2] = -3;
        layer_2_biases[3] = -2;
        layer_2_biases[4] = 8;
        layer_2_biases[5] = 12;
        layer_2_biases[6] = -1;
        layer_2_biases[7] = 0;
        layer_2_biases[8] = -21;
        layer_2_biases[9] = 0;
    end

    integer i, j, k;
    always @(*) begin
        if (predict) begin

            // Layer 1 Computation
            for (j = 0; j < 16; j = j + 1) begin
                layer_1_outputs[j] = layer_1_biases[j]; // Initialize with bias
                for (k = 0; k < 144; k = k + 1) begin
                    if (inp[k] == 1)
                        layer_1_outputs[j] = layer_1_outputs[j] + layer_1_weights[k][j];
                end
            end

            // Layer 2 Computation
            for (j = 0; j < 10; j = j + 1) begin
                layer_2_outputs[j] = layer_2_biases[j]; // Initialize with bias
                for (k = 0; k < 16; k = k + 1) begin
                    layer_2_outputs[j] = layer_2_outputs[j] + layer_1_outputs[k] * layer_2_weights[k][j];
                end
                // Apply ReLU
                if (layer_2_outputs[j] < 0)
                    layer_2_outputs[j] = 0;
            end

            // Winner-takes-all logic
            max_val = layer_2_outputs[0];
            max_idx = 0;
            for (i = 1; i < 10; i = i + 1) begin
                if (layer_2_outputs[i] > max_val) begin
                    max_val = layer_2_outputs[i];
                    max_idx = i;
                end
            end
            class = max_idx;

        end else begin
            class = 10;
        end
    end

endmodule
