module MLP_model (
    input wire [143:0] inp,
    output wire [3:0] class
);

    // Layer 1: Dense
    wire signed [5:0] layer_1_weights [31:0][143:0];
    wire signed [5:0] layer_1_biases [31:0];

    assign layer_1_weights[0][0] = -6'sd1;
    assign layer_1_weights[0][1] = 6'sd1;
    assign layer_1_weights[0][2] = -6'sd1;
    assign layer_1_weights[0][3] = -6'sd7;
    assign layer_1_weights[0][4] = -6'sd5;
    assign layer_1_weights[0][5] = -6'sd3;
    assign layer_1_weights[0][6] = 6'sd0;
    assign layer_1_weights[0][7] = -6'sd2;
    assign layer_1_weights[0][8] = 6'sd1;
    assign layer_1_weights[0][9] = -6'sd8;
    assign layer_1_weights[0][10] = 6'sd0;
    assign layer_1_weights[0][11] = 6'sd0;
    assign layer_1_weights[0][12] = 6'sd0;
    assign layer_1_weights[0][13] = 6'sd2;
    assign layer_1_weights[0][14] = -6'sd4;
    assign layer_1_weights[0][15] = -6'sd3;
    assign layer_1_weights[0][16] = 6'sd1;
    assign layer_1_weights[0][17] = 6'sd0;
    assign layer_1_weights[0][18] = 6'sd0;
    assign layer_1_weights[0][19] = 6'sd5;
    assign layer_1_weights[0][20] = 6'sd2;
    assign layer_1_weights[0][21] = -6'sd2;
    assign layer_1_weights[0][22] = -6'sd2;
    assign layer_1_weights[0][23] = -6'sd1;
    assign layer_1_weights[0][24] = -6'sd1;
    assign layer_1_weights[0][25] = 6'sd0;
    assign layer_1_weights[0][26] = -6'sd5;
    assign layer_1_weights[0][27] = -6'sd1;
    assign layer_1_weights[0][28] = -6'sd1;
    assign layer_1_weights[0][29] = -6'sd2;
    assign layer_1_weights[0][30] = -6'sd1;
    assign layer_1_weights[0][31] = 6'sd0;
    assign layer_1_weights[0][32] = 6'sd4;
    assign layer_1_weights[0][33] = 6'sd3;
    assign layer_1_weights[0][34] = 6'sd3;
    assign layer_1_weights[0][35] = -6'sd8;
    assign layer_1_weights[0][36] = -6'sd5;
    assign layer_1_weights[0][37] = 6'sd4;
    assign layer_1_weights[0][38] = 6'sd0;
    assign layer_1_weights[0][39] = -6'sd1;
    assign layer_1_weights[0][40] = -6'sd1;
    assign layer_1_weights[0][41] = -6'sd3;
    assign layer_1_weights[0][42] = -6'sd7;
    assign layer_1_weights[0][43] = 6'sd4;
    assign layer_1_weights[0][44] = 6'sd6;
    assign layer_1_weights[0][45] = -6'sd1;
    assign layer_1_weights[0][46] = 6'sd4;
    assign layer_1_weights[0][47] = -6'sd1;
    assign layer_1_weights[0][48] = 6'sd4;
    assign layer_1_weights[0][49] = -6'sd4;
    assign layer_1_weights[0][50] = -6'sd2;
    assign layer_1_weights[0][51] = -6'sd2;
    assign layer_1_weights[0][52] = -6'sd1;
    assign layer_1_weights[0][53] = -6'sd6;
    assign layer_1_weights[0][54] = -6'sd5;
    assign layer_1_weights[0][55] = 6'sd6;
    assign layer_1_weights[0][56] = 6'sd4;
    assign layer_1_weights[0][57] = -6'sd2;
    assign layer_1_weights[0][58] = -6'sd4;
    assign layer_1_weights[0][59] = -6'sd3;
    assign layer_1_weights[0][60] = -6'sd1;
    assign layer_1_weights[0][61] = 6'sd0;
    assign layer_1_weights[0][62] = -6'sd2;
    assign layer_1_weights[0][63] = -6'sd2;
    assign layer_1_weights[0][64] = -6'sd5;
    assign layer_1_weights[0][65] = -6'sd4;
    assign layer_1_weights[0][66] = -6'sd7;
    assign layer_1_weights[0][67] = -6'sd1;
    assign layer_1_weights[0][68] = 6'sd0;
    assign layer_1_weights[0][69] = -6'sd1;
    assign layer_1_weights[0][70] = -6'sd4;
    assign layer_1_weights[0][71] = 6'sd0;
    assign layer_1_weights[0][72] = 6'sd2;
    assign layer_1_weights[0][73] = 6'sd2;
    assign layer_1_weights[0][74] = 6'sd4;
    assign layer_1_weights[0][75] = 6'sd1;
    assign layer_1_weights[0][76] = 6'sd0;
    assign layer_1_weights[0][77] = 6'sd2;
    assign layer_1_weights[0][78] = -6'sd2;
    assign layer_1_weights[0][79] = 6'sd1;
    assign layer_1_weights[0][80] = 6'sd2;
    assign layer_1_weights[0][81] = 6'sd0;
    assign layer_1_weights[0][82] = 6'sd0;
    assign layer_1_weights[0][83] = -6'sd2;
    assign layer_1_weights[0][84] = 6'sd5;
    assign layer_1_weights[0][85] = 6'sd3;
    assign layer_1_weights[0][86] = 6'sd8;
    assign layer_1_weights[0][87] = 6'sd6;
    assign layer_1_weights[0][88] = 6'sd4;
    assign layer_1_weights[0][89] = 6'sd9;
    assign layer_1_weights[0][90] = 6'sd2;
    assign layer_1_weights[0][91] = 6'sd0;
    assign layer_1_weights[0][92] = 6'sd0;
    assign layer_1_weights[0][93] = -6'sd2;
    assign layer_1_weights[0][94] = -6'sd5;
    assign layer_1_weights[0][95] = 6'sd7;
    assign layer_1_weights[0][96] = -6'sd2;
    assign layer_1_weights[0][97] = 6'sd1;
    assign layer_1_weights[0][98] = 6'sd4;
    assign layer_1_weights[0][99] = 6'sd1;
    assign layer_1_weights[0][100] = -6'sd1;
    assign layer_1_weights[0][101] = 6'sd2;
    assign layer_1_weights[0][102] = -6'sd3;
    assign layer_1_weights[0][103] = 6'sd2;
    assign layer_1_weights[0][104] = 6'sd3;
    assign layer_1_weights[0][105] = -6'sd4;
    assign layer_1_weights[0][106] = -6'sd1;
    assign layer_1_weights[0][107] = 6'sd4;
    assign layer_1_weights[0][108] = 6'sd7;
    assign layer_1_weights[0][109] = 6'sd0;
    assign layer_1_weights[0][110] = -6'sd1;
    assign layer_1_weights[0][111] = -6'sd2;
    assign layer_1_weights[0][112] = -6'sd1;
    assign layer_1_weights[0][113] = -6'sd1;
    assign layer_1_weights[0][114] = 6'sd0;
    assign layer_1_weights[0][115] = 6'sd3;
    assign layer_1_weights[0][116] = 6'sd4;
    assign layer_1_weights[0][117] = 6'sd8;
    assign layer_1_weights[0][118] = 6'sd4;
    assign layer_1_weights[0][119] = 6'sd4;
    assign layer_1_weights[0][120] = 6'sd0;
    assign layer_1_weights[0][121] = 6'sd2;
    assign layer_1_weights[0][122] = -6'sd2;
    assign layer_1_weights[0][123] = 6'sd0;
    assign layer_1_weights[0][124] = 6'sd2;
    assign layer_1_weights[0][125] = 6'sd1;
    assign layer_1_weights[0][126] = -6'sd1;
    assign layer_1_weights[0][127] = -6'sd1;
    assign layer_1_weights[0][128] = 6'sd0;
    assign layer_1_weights[0][129] = 6'sd2;
    assign layer_1_weights[0][130] = 6'sd3;
    assign layer_1_weights[0][131] = 6'sd7;
    assign layer_1_weights[0][132] = 6'sd1;
    assign layer_1_weights[0][133] = -6'sd1;
    assign layer_1_weights[0][134] = -6'sd4;
    assign layer_1_weights[0][135] = 6'sd4;
    assign layer_1_weights[0][136] = 6'sd1;
    assign layer_1_weights[0][137] = 6'sd7;
    assign layer_1_weights[0][138] = 6'sd4;
    assign layer_1_weights[0][139] = -6'sd4;
    assign layer_1_weights[0][140] = -6'sd2;
    assign layer_1_weights[0][141] = 6'sd1;
    assign layer_1_weights[0][142] = -6'sd1;
    assign layer_1_weights[0][143] = -6'sd1;
    assign layer_1_biases[0] = 6'sd3;
    assign layer_1_weights[1][0] = 6'sd0;
    assign layer_1_weights[1][1] = 6'sd0;
    assign layer_1_weights[1][2] = 6'sd0;
    assign layer_1_weights[1][3] = -6'sd3;
    assign layer_1_weights[1][4] = 6'sd2;
    assign layer_1_weights[1][5] = -6'sd4;
    assign layer_1_weights[1][6] = 6'sd4;
    assign layer_1_weights[1][7] = -6'sd2;
    assign layer_1_weights[1][8] = 6'sd7;
    assign layer_1_weights[1][9] = -6'sd2;
    assign layer_1_weights[1][10] = -6'sd1;
    assign layer_1_weights[1][11] = -6'sd2;
    assign layer_1_weights[1][12] = 6'sd0;
    assign layer_1_weights[1][13] = -6'sd1;
    assign layer_1_weights[1][14] = 6'sd4;
    assign layer_1_weights[1][15] = 6'sd4;
    assign layer_1_weights[1][16] = 6'sd6;
    assign layer_1_weights[1][17] = 6'sd6;
    assign layer_1_weights[1][18] = 6'sd5;
    assign layer_1_weights[1][19] = 6'sd1;
    assign layer_1_weights[1][20] = 6'sd3;
    assign layer_1_weights[1][21] = 6'sd4;
    assign layer_1_weights[1][22] = 6'sd2;
    assign layer_1_weights[1][23] = 6'sd1;
    assign layer_1_weights[1][24] = -6'sd1;
    assign layer_1_weights[1][25] = -6'sd4;
    assign layer_1_weights[1][26] = 6'sd2;
    assign layer_1_weights[1][27] = 6'sd0;
    assign layer_1_weights[1][28] = 6'sd4;
    assign layer_1_weights[1][29] = 6'sd3;
    assign layer_1_weights[1][30] = 6'sd2;
    assign layer_1_weights[1][31] = 6'sd3;
    assign layer_1_weights[1][32] = 6'sd1;
    assign layer_1_weights[1][33] = 6'sd1;
    assign layer_1_weights[1][34] = 6'sd3;
    assign layer_1_weights[1][35] = 6'sd7;
    assign layer_1_weights[1][36] = 6'sd2;
    assign layer_1_weights[1][37] = -6'sd2;
    assign layer_1_weights[1][38] = 6'sd1;
    assign layer_1_weights[1][39] = 6'sd0;
    assign layer_1_weights[1][40] = 6'sd1;
    assign layer_1_weights[1][41] = 6'sd0;
    assign layer_1_weights[1][42] = 6'sd0;
    assign layer_1_weights[1][43] = -6'sd1;
    assign layer_1_weights[1][44] = -6'sd1;
    assign layer_1_weights[1][45] = 6'sd1;
    assign layer_1_weights[1][46] = 6'sd1;
    assign layer_1_weights[1][47] = 6'sd6;
    assign layer_1_weights[1][48] = -6'sd3;
    assign layer_1_weights[1][49] = 6'sd4;
    assign layer_1_weights[1][50] = 6'sd1;
    assign layer_1_weights[1][51] = 6'sd0;
    assign layer_1_weights[1][52] = -6'sd3;
    assign layer_1_weights[1][53] = -6'sd1;
    assign layer_1_weights[1][54] = 6'sd1;
    assign layer_1_weights[1][55] = -6'sd1;
    assign layer_1_weights[1][56] = -6'sd3;
    assign layer_1_weights[1][57] = -6'sd1;
    assign layer_1_weights[1][58] = -6'sd1;
    assign layer_1_weights[1][59] = -6'sd6;
    assign layer_1_weights[1][60] = -6'sd6;
    assign layer_1_weights[1][61] = -6'sd2;
    assign layer_1_weights[1][62] = -6'sd2;
    assign layer_1_weights[1][63] = 6'sd0;
    assign layer_1_weights[1][64] = 6'sd3;
    assign layer_1_weights[1][65] = 6'sd4;
    assign layer_1_weights[1][66] = 6'sd4;
    assign layer_1_weights[1][67] = 6'sd0;
    assign layer_1_weights[1][68] = 6'sd1;
    assign layer_1_weights[1][69] = 6'sd2;
    assign layer_1_weights[1][70] = -6'sd6;
    assign layer_1_weights[1][71] = -6'sd10;
    assign layer_1_weights[1][72] = 6'sd4;
    assign layer_1_weights[1][73] = 6'sd1;
    assign layer_1_weights[1][74] = -6'sd4;
    assign layer_1_weights[1][75] = -6'sd9;
    assign layer_1_weights[1][76] = -6'sd7;
    assign layer_1_weights[1][77] = -6'sd6;
    assign layer_1_weights[1][78] = -6'sd2;
    assign layer_1_weights[1][79] = -6'sd4;
    assign layer_1_weights[1][80] = 6'sd2;
    assign layer_1_weights[1][81] = 6'sd3;
    assign layer_1_weights[1][82] = -6'sd1;
    assign layer_1_weights[1][83] = -6'sd4;
    assign layer_1_weights[1][84] = 6'sd7;
    assign layer_1_weights[1][85] = 6'sd0;
    assign layer_1_weights[1][86] = -6'sd2;
    assign layer_1_weights[1][87] = -6'sd8;
    assign layer_1_weights[1][88] = -6'sd13;
    assign layer_1_weights[1][89] = -6'sd9;
    assign layer_1_weights[1][90] = -6'sd4;
    assign layer_1_weights[1][91] = 6'sd0;
    assign layer_1_weights[1][92] = 6'sd0;
    assign layer_1_weights[1][93] = 6'sd0;
    assign layer_1_weights[1][94] = 6'sd0;
    assign layer_1_weights[1][95] = 6'sd4;
    assign layer_1_weights[1][96] = 6'sd4;
    assign layer_1_weights[1][97] = 6'sd3;
    assign layer_1_weights[1][98] = 6'sd6;
    assign layer_1_weights[1][99] = 6'sd7;
    assign layer_1_weights[1][100] = 6'sd3;
    assign layer_1_weights[1][101] = 6'sd6;
    assign layer_1_weights[1][102] = 6'sd4;
    assign layer_1_weights[1][103] = 6'sd2;
    assign layer_1_weights[1][104] = -6'sd1;
    assign layer_1_weights[1][105] = 6'sd0;
    assign layer_1_weights[1][106] = 6'sd3;
    assign layer_1_weights[1][107] = 6'sd3;
    assign layer_1_weights[1][108] = -6'sd3;
    assign layer_1_weights[1][109] = 6'sd5;
    assign layer_1_weights[1][110] = 6'sd4;
    assign layer_1_weights[1][111] = 6'sd5;
    assign layer_1_weights[1][112] = 6'sd7;
    assign layer_1_weights[1][113] = 6'sd2;
    assign layer_1_weights[1][114] = 6'sd0;
    assign layer_1_weights[1][115] = 6'sd2;
    assign layer_1_weights[1][116] = 6'sd0;
    assign layer_1_weights[1][117] = -6'sd1;
    assign layer_1_weights[1][118] = 6'sd5;
    assign layer_1_weights[1][119] = -6'sd8;
    assign layer_1_weights[1][120] = 6'sd1;
    assign layer_1_weights[1][121] = 6'sd4;
    assign layer_1_weights[1][122] = -6'sd7;
    assign layer_1_weights[1][123] = -6'sd3;
    assign layer_1_weights[1][124] = -6'sd2;
    assign layer_1_weights[1][125] = -6'sd1;
    assign layer_1_weights[1][126] = -6'sd1;
    assign layer_1_weights[1][127] = 6'sd2;
    assign layer_1_weights[1][128] = 6'sd2;
    assign layer_1_weights[1][129] = -6'sd1;
    assign layer_1_weights[1][130] = 6'sd5;
    assign layer_1_weights[1][131] = 6'sd0;
    assign layer_1_weights[1][132] = 6'sd1;
    assign layer_1_weights[1][133] = -6'sd1;
    assign layer_1_weights[1][134] = -6'sd1;
    assign layer_1_weights[1][135] = 6'sd0;
    assign layer_1_weights[1][136] = 6'sd2;
    assign layer_1_weights[1][137] = 6'sd3;
    assign layer_1_weights[1][138] = 6'sd2;
    assign layer_1_weights[1][139] = -6'sd1;
    assign layer_1_weights[1][140] = -6'sd3;
    assign layer_1_weights[1][141] = -6'sd5;
    assign layer_1_weights[1][142] = 6'sd2;
    assign layer_1_weights[1][143] = 6'sd2;
    assign layer_1_biases[1] = -6'sd1;
    assign layer_1_weights[2][0] = -6'sd1;
    assign layer_1_weights[2][1] = 6'sd0;
    assign layer_1_weights[2][2] = -6'sd1;
    assign layer_1_weights[2][3] = -6'sd1;
    assign layer_1_weights[2][4] = 6'sd2;
    assign layer_1_weights[2][5] = 6'sd7;
    assign layer_1_weights[2][6] = 6'sd3;
    assign layer_1_weights[2][7] = -6'sd3;
    assign layer_1_weights[2][8] = -6'sd2;
    assign layer_1_weights[2][9] = 6'sd0;
    assign layer_1_weights[2][10] = 6'sd1;
    assign layer_1_weights[2][11] = -6'sd1;
    assign layer_1_weights[2][12] = 6'sd2;
    assign layer_1_weights[2][13] = -6'sd2;
    assign layer_1_weights[2][14] = 6'sd5;
    assign layer_1_weights[2][15] = 6'sd6;
    assign layer_1_weights[2][16] = 6'sd0;
    assign layer_1_weights[2][17] = -6'sd1;
    assign layer_1_weights[2][18] = -6'sd2;
    assign layer_1_weights[2][19] = -6'sd2;
    assign layer_1_weights[2][20] = 6'sd1;
    assign layer_1_weights[2][21] = -6'sd4;
    assign layer_1_weights[2][22] = -6'sd3;
    assign layer_1_weights[2][23] = -6'sd3;
    assign layer_1_weights[2][24] = 6'sd0;
    assign layer_1_weights[2][25] = 6'sd0;
    assign layer_1_weights[2][26] = 6'sd1;
    assign layer_1_weights[2][27] = 6'sd0;
    assign layer_1_weights[2][28] = 6'sd0;
    assign layer_1_weights[2][29] = 6'sd1;
    assign layer_1_weights[2][30] = -6'sd1;
    assign layer_1_weights[2][31] = 6'sd2;
    assign layer_1_weights[2][32] = -6'sd1;
    assign layer_1_weights[2][33] = -6'sd4;
    assign layer_1_weights[2][34] = 6'sd1;
    assign layer_1_weights[2][35] = -6'sd7;
    assign layer_1_weights[2][36] = 6'sd0;
    assign layer_1_weights[2][37] = 6'sd6;
    assign layer_1_weights[2][38] = 6'sd2;
    assign layer_1_weights[2][39] = 6'sd2;
    assign layer_1_weights[2][40] = 6'sd4;
    assign layer_1_weights[2][41] = -6'sd1;
    assign layer_1_weights[2][42] = 6'sd0;
    assign layer_1_weights[2][43] = 6'sd5;
    assign layer_1_weights[2][44] = 6'sd1;
    assign layer_1_weights[2][45] = -6'sd1;
    assign layer_1_weights[2][46] = -6'sd4;
    assign layer_1_weights[2][47] = 6'sd0;
    assign layer_1_weights[2][48] = 6'sd6;
    assign layer_1_weights[2][49] = 6'sd2;
    assign layer_1_weights[2][50] = -6'sd1;
    assign layer_1_weights[2][51] = 6'sd4;
    assign layer_1_weights[2][52] = -6'sd4;
    assign layer_1_weights[2][53] = -6'sd3;
    assign layer_1_weights[2][54] = 6'sd2;
    assign layer_1_weights[2][55] = 6'sd2;
    assign layer_1_weights[2][56] = -6'sd2;
    assign layer_1_weights[2][57] = -6'sd1;
    assign layer_1_weights[2][58] = -6'sd2;
    assign layer_1_weights[2][59] = -6'sd1;
    assign layer_1_weights[2][60] = -6'sd2;
    assign layer_1_weights[2][61] = -6'sd3;
    assign layer_1_weights[2][62] = 6'sd3;
    assign layer_1_weights[2][63] = -6'sd4;
    assign layer_1_weights[2][64] = -6'sd1;
    assign layer_1_weights[2][65] = 6'sd2;
    assign layer_1_weights[2][66] = 6'sd8;
    assign layer_1_weights[2][67] = 6'sd1;
    assign layer_1_weights[2][68] = 6'sd0;
    assign layer_1_weights[2][69] = -6'sd1;
    assign layer_1_weights[2][70] = 6'sd0;
    assign layer_1_weights[2][71] = -6'sd4;
    assign layer_1_weights[2][72] = 6'sd1;
    assign layer_1_weights[2][73] = -6'sd1;
    assign layer_1_weights[2][74] = -6'sd3;
    assign layer_1_weights[2][75] = 6'sd3;
    assign layer_1_weights[2][76] = 6'sd8;
    assign layer_1_weights[2][77] = 6'sd8;
    assign layer_1_weights[2][78] = 6'sd4;
    assign layer_1_weights[2][79] = 6'sd3;
    assign layer_1_weights[2][80] = 6'sd0;
    assign layer_1_weights[2][81] = 6'sd1;
    assign layer_1_weights[2][82] = -6'sd7;
    assign layer_1_weights[2][83] = -6'sd5;
    assign layer_1_weights[2][84] = 6'sd2;
    assign layer_1_weights[2][85] = -6'sd10;
    assign layer_1_weights[2][86] = -6'sd15;
    assign layer_1_weights[2][87] = -6'sd13;
    assign layer_1_weights[2][88] = -6'sd5;
    assign layer_1_weights[2][89] = -6'sd1;
    assign layer_1_weights[2][90] = 6'sd2;
    assign layer_1_weights[2][91] = -6'sd2;
    assign layer_1_weights[2][92] = -6'sd5;
    assign layer_1_weights[2][93] = -6'sd1;
    assign layer_1_weights[2][94] = -6'sd2;
    assign layer_1_weights[2][95] = -6'sd3;
    assign layer_1_weights[2][96] = 6'sd9;
    assign layer_1_weights[2][97] = 6'sd3;
    assign layer_1_weights[2][98] = -6'sd1;
    assign layer_1_weights[2][99] = -6'sd5;
    assign layer_1_weights[2][100] = -6'sd8;
    assign layer_1_weights[2][101] = -6'sd7;
    assign layer_1_weights[2][102] = -6'sd2;
    assign layer_1_weights[2][103] = -6'sd3;
    assign layer_1_weights[2][104] = -6'sd3;
    assign layer_1_weights[2][105] = -6'sd1;
    assign layer_1_weights[2][106] = -6'sd3;
    assign layer_1_weights[2][107] = 6'sd5;
    assign layer_1_weights[2][108] = 6'sd2;
    assign layer_1_weights[2][109] = 6'sd7;
    assign layer_1_weights[2][110] = 6'sd5;
    assign layer_1_weights[2][111] = 6'sd3;
    assign layer_1_weights[2][112] = 6'sd1;
    assign layer_1_weights[2][113] = -6'sd2;
    assign layer_1_weights[2][114] = -6'sd1;
    assign layer_1_weights[2][115] = -6'sd3;
    assign layer_1_weights[2][116] = -6'sd2;
    assign layer_1_weights[2][117] = -6'sd2;
    assign layer_1_weights[2][118] = -6'sd4;
    assign layer_1_weights[2][119] = 6'sd6;
    assign layer_1_weights[2][120] = -6'sd1;
    assign layer_1_weights[2][121] = 6'sd9;
    assign layer_1_weights[2][122] = 6'sd4;
    assign layer_1_weights[2][123] = 6'sd3;
    assign layer_1_weights[2][124] = 6'sd1;
    assign layer_1_weights[2][125] = 6'sd0;
    assign layer_1_weights[2][126] = -6'sd1;
    assign layer_1_weights[2][127] = 6'sd0;
    assign layer_1_weights[2][128] = 6'sd2;
    assign layer_1_weights[2][129] = -6'sd2;
    assign layer_1_weights[2][130] = -6'sd3;
    assign layer_1_weights[2][131] = -6'sd1;
    assign layer_1_weights[2][132] = 6'sd1;
    assign layer_1_weights[2][133] = 6'sd3;
    assign layer_1_weights[2][134] = 6'sd6;
    assign layer_1_weights[2][135] = 6'sd0;
    assign layer_1_weights[2][136] = 6'sd1;
    assign layer_1_weights[2][137] = -6'sd5;
    assign layer_1_weights[2][138] = 6'sd2;
    assign layer_1_weights[2][139] = -6'sd2;
    assign layer_1_weights[2][140] = 6'sd1;
    assign layer_1_weights[2][141] = 6'sd0;
    assign layer_1_weights[2][142] = 6'sd2;
    assign layer_1_weights[2][143] = 6'sd1;
    assign layer_1_biases[2] = 6'sd2;
    assign layer_1_weights[3][0] = 6'sd1;
    assign layer_1_weights[3][1] = 6'sd0;
    assign layer_1_weights[3][2] = -6'sd3;
    assign layer_1_weights[3][3] = -6'sd4;
    assign layer_1_weights[3][4] = -6'sd1;
    assign layer_1_weights[3][5] = -6'sd11;
    assign layer_1_weights[3][6] = 6'sd2;
    assign layer_1_weights[3][7] = 6'sd1;
    assign layer_1_weights[3][8] = -6'sd1;
    assign layer_1_weights[3][9] = -6'sd2;
    assign layer_1_weights[3][10] = -6'sd1;
    assign layer_1_weights[3][11] = 6'sd1;
    assign layer_1_weights[3][12] = 6'sd1;
    assign layer_1_weights[3][13] = 6'sd2;
    assign layer_1_weights[3][14] = 6'sd7;
    assign layer_1_weights[3][15] = 6'sd2;
    assign layer_1_weights[3][16] = 6'sd1;
    assign layer_1_weights[3][17] = 6'sd2;
    assign layer_1_weights[3][18] = -6'sd5;
    assign layer_1_weights[3][19] = -6'sd7;
    assign layer_1_weights[3][20] = -6'sd14;
    assign layer_1_weights[3][21] = -6'sd5;
    assign layer_1_weights[3][22] = -6'sd3;
    assign layer_1_weights[3][23] = 6'sd2;
    assign layer_1_weights[3][24] = 6'sd0;
    assign layer_1_weights[3][25] = 6'sd6;
    assign layer_1_weights[3][26] = 6'sd3;
    assign layer_1_weights[3][27] = 6'sd1;
    assign layer_1_weights[3][28] = 6'sd3;
    assign layer_1_weights[3][29] = 6'sd4;
    assign layer_1_weights[3][30] = 6'sd0;
    assign layer_1_weights[3][31] = -6'sd7;
    assign layer_1_weights[3][32] = -6'sd9;
    assign layer_1_weights[3][33] = -6'sd9;
    assign layer_1_weights[3][34] = -6'sd7;
    assign layer_1_weights[3][35] = -6'sd6;
    assign layer_1_weights[3][36] = 6'sd6;
    assign layer_1_weights[3][37] = 6'sd8;
    assign layer_1_weights[3][38] = 6'sd2;
    assign layer_1_weights[3][39] = 6'sd1;
    assign layer_1_weights[3][40] = 6'sd1;
    assign layer_1_weights[3][41] = 6'sd4;
    assign layer_1_weights[3][42] = 6'sd7;
    assign layer_1_weights[3][43] = 6'sd3;
    assign layer_1_weights[3][44] = -6'sd10;
    assign layer_1_weights[3][45] = -6'sd19;
    assign layer_1_weights[3][46] = -6'sd8;
    assign layer_1_weights[3][47] = -6'sd3;
    assign layer_1_weights[3][48] = 6'sd9;
    assign layer_1_weights[3][49] = 6'sd0;
    assign layer_1_weights[3][50] = 6'sd2;
    assign layer_1_weights[3][51] = -6'sd2;
    assign layer_1_weights[3][52] = -6'sd2;
    assign layer_1_weights[3][53] = 6'sd0;
    assign layer_1_weights[3][54] = 6'sd7;
    assign layer_1_weights[3][55] = 6'sd5;
    assign layer_1_weights[3][56] = -6'sd7;
    assign layer_1_weights[3][57] = -6'sd16;
    assign layer_1_weights[3][58] = 6'sd1;
    assign layer_1_weights[3][59] = 6'sd9;
    assign layer_1_weights[3][60] = 6'sd8;
    assign layer_1_weights[3][61] = 6'sd0;
    assign layer_1_weights[3][62] = -6'sd3;
    assign layer_1_weights[3][63] = 6'sd1;
    assign layer_1_weights[3][64] = -6'sd2;
    assign layer_1_weights[3][65] = -6'sd3;
    assign layer_1_weights[3][66] = 6'sd2;
    assign layer_1_weights[3][67] = 6'sd3;
    assign layer_1_weights[3][68] = -6'sd8;
    assign layer_1_weights[3][69] = -6'sd10;
    assign layer_1_weights[3][70] = 6'sd0;
    assign layer_1_weights[3][71] = 6'sd8;
    assign layer_1_weights[3][72] = 6'sd1;
    assign layer_1_weights[3][73] = -6'sd3;
    assign layer_1_weights[3][74] = -6'sd2;
    assign layer_1_weights[3][75] = 6'sd3;
    assign layer_1_weights[3][76] = -6'sd4;
    assign layer_1_weights[3][77] = -6'sd1;
    assign layer_1_weights[3][78] = 6'sd6;
    assign layer_1_weights[3][79] = 6'sd0;
    assign layer_1_weights[3][80] = -6'sd6;
    assign layer_1_weights[3][81] = 6'sd3;
    assign layer_1_weights[3][82] = 6'sd0;
    assign layer_1_weights[3][83] = 6'sd1;
    assign layer_1_weights[3][84] = 6'sd1;
    assign layer_1_weights[3][85] = -6'sd3;
    assign layer_1_weights[3][86] = 6'sd2;
    assign layer_1_weights[3][87] = -6'sd1;
    assign layer_1_weights[3][88] = -6'sd1;
    assign layer_1_weights[3][89] = -6'sd1;
    assign layer_1_weights[3][90] = 6'sd4;
    assign layer_1_weights[3][91] = 6'sd0;
    assign layer_1_weights[3][92] = 6'sd3;
    assign layer_1_weights[3][93] = 6'sd2;
    assign layer_1_weights[3][94] = 6'sd3;
    assign layer_1_weights[3][95] = 6'sd0;
    assign layer_1_weights[3][96] = 6'sd7;
    assign layer_1_weights[3][97] = -6'sd1;
    assign layer_1_weights[3][98] = 6'sd1;
    assign layer_1_weights[3][99] = -6'sd1;
    assign layer_1_weights[3][100] = -6'sd3;
    assign layer_1_weights[3][101] = -6'sd2;
    assign layer_1_weights[3][102] = 6'sd3;
    assign layer_1_weights[3][103] = -6'sd1;
    assign layer_1_weights[3][104] = 6'sd2;
    assign layer_1_weights[3][105] = 6'sd4;
    assign layer_1_weights[3][106] = 6'sd0;
    assign layer_1_weights[3][107] = 6'sd5;
    assign layer_1_weights[3][108] = 6'sd7;
    assign layer_1_weights[3][109] = 6'sd5;
    assign layer_1_weights[3][110] = -6'sd3;
    assign layer_1_weights[3][111] = 6'sd2;
    assign layer_1_weights[3][112] = 6'sd3;
    assign layer_1_weights[3][113] = 6'sd2;
    assign layer_1_weights[3][114] = -6'sd1;
    assign layer_1_weights[3][115] = 6'sd0;
    assign layer_1_weights[3][116] = 6'sd0;
    assign layer_1_weights[3][117] = 6'sd2;
    assign layer_1_weights[3][118] = -6'sd1;
    assign layer_1_weights[3][119] = -6'sd7;
    assign layer_1_weights[3][120] = 6'sd0;
    assign layer_1_weights[3][121] = 6'sd3;
    assign layer_1_weights[3][122] = -6'sd3;
    assign layer_1_weights[3][123] = 6'sd0;
    assign layer_1_weights[3][124] = 6'sd0;
    assign layer_1_weights[3][125] = 6'sd1;
    assign layer_1_weights[3][126] = 6'sd0;
    assign layer_1_weights[3][127] = 6'sd0;
    assign layer_1_weights[3][128] = 6'sd3;
    assign layer_1_weights[3][129] = 6'sd0;
    assign layer_1_weights[3][130] = 6'sd1;
    assign layer_1_weights[3][131] = 6'sd8;
    assign layer_1_weights[3][132] = 6'sd0;
    assign layer_1_weights[3][133] = 6'sd0;
    assign layer_1_weights[3][134] = 6'sd7;
    assign layer_1_weights[3][135] = 6'sd7;
    assign layer_1_weights[3][136] = 6'sd3;
    assign layer_1_weights[3][137] = -6'sd1;
    assign layer_1_weights[3][138] = -6'sd6;
    assign layer_1_weights[3][139] = -6'sd1;
    assign layer_1_weights[3][140] = 6'sd2;
    assign layer_1_weights[3][141] = -6'sd6;
    assign layer_1_weights[3][142] = 6'sd0;
    assign layer_1_weights[3][143] = -6'sd1;
    assign layer_1_biases[3] = 6'sd5;
    assign layer_1_weights[4][0] = 6'sd0;
    assign layer_1_weights[4][1] = 6'sd0;
    assign layer_1_weights[4][2] = -6'sd4;
    assign layer_1_weights[4][3] = -6'sd7;
    assign layer_1_weights[4][4] = -6'sd11;
    assign layer_1_weights[4][5] = -6'sd6;
    assign layer_1_weights[4][6] = -6'sd6;
    assign layer_1_weights[4][7] = -6'sd5;
    assign layer_1_weights[4][8] = -6'sd2;
    assign layer_1_weights[4][9] = -6'sd5;
    assign layer_1_weights[4][10] = 6'sd1;
    assign layer_1_weights[4][11] = -6'sd1;
    assign layer_1_weights[4][12] = 6'sd0;
    assign layer_1_weights[4][13] = 6'sd0;
    assign layer_1_weights[4][14] = -6'sd2;
    assign layer_1_weights[4][15] = -6'sd3;
    assign layer_1_weights[4][16] = 6'sd1;
    assign layer_1_weights[4][17] = -6'sd3;
    assign layer_1_weights[4][18] = -6'sd4;
    assign layer_1_weights[4][19] = 6'sd1;
    assign layer_1_weights[4][20] = -6'sd1;
    assign layer_1_weights[4][21] = -6'sd1;
    assign layer_1_weights[4][22] = 6'sd3;
    assign layer_1_weights[4][23] = -6'sd4;
    assign layer_1_weights[4][24] = -6'sd1;
    assign layer_1_weights[4][25] = -6'sd5;
    assign layer_1_weights[4][26] = 6'sd2;
    assign layer_1_weights[4][27] = -6'sd2;
    assign layer_1_weights[4][28] = 6'sd0;
    assign layer_1_weights[4][29] = 6'sd0;
    assign layer_1_weights[4][30] = -6'sd2;
    assign layer_1_weights[4][31] = 6'sd0;
    assign layer_1_weights[4][32] = 6'sd3;
    assign layer_1_weights[4][33] = -6'sd1;
    assign layer_1_weights[4][34] = 6'sd1;
    assign layer_1_weights[4][35] = -6'sd8;
    assign layer_1_weights[4][36] = 6'sd3;
    assign layer_1_weights[4][37] = 6'sd4;
    assign layer_1_weights[4][38] = 6'sd1;
    assign layer_1_weights[4][39] = 6'sd2;
    assign layer_1_weights[4][40] = 6'sd0;
    assign layer_1_weights[4][41] = -6'sd3;
    assign layer_1_weights[4][42] = -6'sd4;
    assign layer_1_weights[4][43] = 6'sd1;
    assign layer_1_weights[4][44] = 6'sd3;
    assign layer_1_weights[4][45] = 6'sd2;
    assign layer_1_weights[4][46] = -6'sd1;
    assign layer_1_weights[4][47] = 6'sd1;
    assign layer_1_weights[4][48] = -6'sd1;
    assign layer_1_weights[4][49] = 6'sd0;
    assign layer_1_weights[4][50] = 6'sd2;
    assign layer_1_weights[4][51] = 6'sd3;
    assign layer_1_weights[4][52] = 6'sd1;
    assign layer_1_weights[4][53] = -6'sd3;
    assign layer_1_weights[4][54] = -6'sd1;
    assign layer_1_weights[4][55] = 6'sd2;
    assign layer_1_weights[4][56] = -6'sd4;
    assign layer_1_weights[4][57] = -6'sd3;
    assign layer_1_weights[4][58] = -6'sd2;
    assign layer_1_weights[4][59] = -6'sd1;
    assign layer_1_weights[4][60] = 6'sd11;
    assign layer_1_weights[4][61] = -6'sd1;
    assign layer_1_weights[4][62] = 6'sd4;
    assign layer_1_weights[4][63] = 6'sd4;
    assign layer_1_weights[4][64] = 6'sd6;
    assign layer_1_weights[4][65] = 6'sd0;
    assign layer_1_weights[4][66] = -6'sd2;
    assign layer_1_weights[4][67] = 6'sd1;
    assign layer_1_weights[4][68] = 6'sd1;
    assign layer_1_weights[4][69] = 6'sd2;
    assign layer_1_weights[4][70] = -6'sd3;
    assign layer_1_weights[4][71] = 6'sd0;
    assign layer_1_weights[4][72] = 6'sd4;
    assign layer_1_weights[4][73] = 6'sd4;
    assign layer_1_weights[4][74] = 6'sd4;
    assign layer_1_weights[4][75] = 6'sd1;
    assign layer_1_weights[4][76] = -6'sd2;
    assign layer_1_weights[4][77] = -6'sd7;
    assign layer_1_weights[4][78] = -6'sd1;
    assign layer_1_weights[4][79] = 6'sd2;
    assign layer_1_weights[4][80] = 6'sd2;
    assign layer_1_weights[4][81] = 6'sd3;
    assign layer_1_weights[4][82] = 6'sd8;
    assign layer_1_weights[4][83] = 6'sd0;
    assign layer_1_weights[4][84] = 6'sd0;
    assign layer_1_weights[4][85] = 6'sd3;
    assign layer_1_weights[4][86] = -6'sd4;
    assign layer_1_weights[4][87] = -6'sd5;
    assign layer_1_weights[4][88] = -6'sd11;
    assign layer_1_weights[4][89] = 6'sd0;
    assign layer_1_weights[4][90] = 6'sd5;
    assign layer_1_weights[4][91] = 6'sd3;
    assign layer_1_weights[4][92] = -6'sd2;
    assign layer_1_weights[4][93] = -6'sd4;
    assign layer_1_weights[4][94] = -6'sd10;
    assign layer_1_weights[4][95] = -6'sd2;
    assign layer_1_weights[4][96] = -6'sd2;
    assign layer_1_weights[4][97] = -6'sd4;
    assign layer_1_weights[4][98] = -6'sd11;
    assign layer_1_weights[4][99] = -6'sd6;
    assign layer_1_weights[4][100] = -6'sd3;
    assign layer_1_weights[4][101] = 6'sd5;
    assign layer_1_weights[4][102] = 6'sd2;
    assign layer_1_weights[4][103] = 6'sd2;
    assign layer_1_weights[4][104] = -6'sd3;
    assign layer_1_weights[4][105] = -6'sd6;
    assign layer_1_weights[4][106] = -6'sd7;
    assign layer_1_weights[4][107] = -6'sd8;
    assign layer_1_weights[4][108] = -6'sd3;
    assign layer_1_weights[4][109] = -6'sd9;
    assign layer_1_weights[4][110] = -6'sd5;
    assign layer_1_weights[4][111] = -6'sd1;
    assign layer_1_weights[4][112] = -6'sd3;
    assign layer_1_weights[4][113] = 6'sd4;
    assign layer_1_weights[4][114] = 6'sd1;
    assign layer_1_weights[4][115] = 6'sd3;
    assign layer_1_weights[4][116] = -6'sd1;
    assign layer_1_weights[4][117] = 6'sd2;
    assign layer_1_weights[4][118] = -6'sd1;
    assign layer_1_weights[4][119] = 6'sd0;
    assign layer_1_weights[4][120] = 6'sd1;
    assign layer_1_weights[4][121] = -6'sd6;
    assign layer_1_weights[4][122] = -6'sd5;
    assign layer_1_weights[4][123] = 6'sd0;
    assign layer_1_weights[4][124] = -6'sd2;
    assign layer_1_weights[4][125] = -6'sd4;
    assign layer_1_weights[4][126] = 6'sd3;
    assign layer_1_weights[4][127] = 6'sd4;
    assign layer_1_weights[4][128] = 6'sd5;
    assign layer_1_weights[4][129] = 6'sd5;
    assign layer_1_weights[4][130] = 6'sd4;
    assign layer_1_weights[4][131] = 6'sd0;
    assign layer_1_weights[4][132] = -6'sd2;
    assign layer_1_weights[4][133] = 6'sd4;
    assign layer_1_weights[4][134] = -6'sd6;
    assign layer_1_weights[4][135] = -6'sd1;
    assign layer_1_weights[4][136] = -6'sd2;
    assign layer_1_weights[4][137] = -6'sd2;
    assign layer_1_weights[4][138] = 6'sd2;
    assign layer_1_weights[4][139] = 6'sd1;
    assign layer_1_weights[4][140] = 6'sd2;
    assign layer_1_weights[4][141] = 6'sd0;
    assign layer_1_weights[4][142] = -6'sd1;
    assign layer_1_weights[4][143] = -6'sd1;
    assign layer_1_biases[4] = 6'sd3;
    assign layer_1_weights[5][0] = 6'sd0;
    assign layer_1_weights[5][1] = -6'sd1;
    assign layer_1_weights[5][2] = -6'sd4;
    assign layer_1_weights[5][3] = -6'sd5;
    assign layer_1_weights[5][4] = -6'sd4;
    assign layer_1_weights[5][5] = 6'sd1;
    assign layer_1_weights[5][6] = -6'sd3;
    assign layer_1_weights[5][7] = -6'sd4;
    assign layer_1_weights[5][8] = -6'sd7;
    assign layer_1_weights[5][9] = -6'sd9;
    assign layer_1_weights[5][10] = -6'sd1;
    assign layer_1_weights[5][11] = 6'sd0;
    assign layer_1_weights[5][12] = -6'sd1;
    assign layer_1_weights[5][13] = 6'sd0;
    assign layer_1_weights[5][14] = -6'sd7;
    assign layer_1_weights[5][15] = -6'sd5;
    assign layer_1_weights[5][16] = 6'sd0;
    assign layer_1_weights[5][17] = -6'sd5;
    assign layer_1_weights[5][18] = -6'sd3;
    assign layer_1_weights[5][19] = 6'sd0;
    assign layer_1_weights[5][20] = -6'sd4;
    assign layer_1_weights[5][21] = -6'sd1;
    assign layer_1_weights[5][22] = -6'sd2;
    assign layer_1_weights[5][23] = 6'sd2;
    assign layer_1_weights[5][24] = 6'sd0;
    assign layer_1_weights[5][25] = 6'sd8;
    assign layer_1_weights[5][26] = -6'sd1;
    assign layer_1_weights[5][27] = 6'sd5;
    assign layer_1_weights[5][28] = -6'sd2;
    assign layer_1_weights[5][29] = -6'sd5;
    assign layer_1_weights[5][30] = 6'sd0;
    assign layer_1_weights[5][31] = 6'sd0;
    assign layer_1_weights[5][32] = -6'sd1;
    assign layer_1_weights[5][33] = -6'sd1;
    assign layer_1_weights[5][34] = -6'sd7;
    assign layer_1_weights[5][35] = 6'sd0;
    assign layer_1_weights[5][36] = 6'sd1;
    assign layer_1_weights[5][37] = 6'sd0;
    assign layer_1_weights[5][38] = 6'sd0;
    assign layer_1_weights[5][39] = 6'sd3;
    assign layer_1_weights[5][40] = -6'sd1;
    assign layer_1_weights[5][41] = -6'sd2;
    assign layer_1_weights[5][42] = 6'sd2;
    assign layer_1_weights[5][43] = 6'sd1;
    assign layer_1_weights[5][44] = -6'sd1;
    assign layer_1_weights[5][45] = -6'sd3;
    assign layer_1_weights[5][46] = -6'sd3;
    assign layer_1_weights[5][47] = -6'sd2;
    assign layer_1_weights[5][48] = -6'sd2;
    assign layer_1_weights[5][49] = -6'sd7;
    assign layer_1_weights[5][50] = 6'sd2;
    assign layer_1_weights[5][51] = 6'sd1;
    assign layer_1_weights[5][52] = 6'sd1;
    assign layer_1_weights[5][53] = 6'sd3;
    assign layer_1_weights[5][54] = 6'sd0;
    assign layer_1_weights[5][55] = 6'sd2;
    assign layer_1_weights[5][56] = 6'sd3;
    assign layer_1_weights[5][57] = -6'sd3;
    assign layer_1_weights[5][58] = -6'sd8;
    assign layer_1_weights[5][59] = -6'sd3;
    assign layer_1_weights[5][60] = 6'sd6;
    assign layer_1_weights[5][61] = 6'sd1;
    assign layer_1_weights[5][62] = 6'sd1;
    assign layer_1_weights[5][63] = 6'sd2;
    assign layer_1_weights[5][64] = 6'sd3;
    assign layer_1_weights[5][65] = 6'sd0;
    assign layer_1_weights[5][66] = 6'sd1;
    assign layer_1_weights[5][67] = 6'sd4;
    assign layer_1_weights[5][68] = 6'sd4;
    assign layer_1_weights[5][69] = -6'sd1;
    assign layer_1_weights[5][70] = -6'sd7;
    assign layer_1_weights[5][71] = -6'sd4;
    assign layer_1_weights[5][72] = 6'sd3;
    assign layer_1_weights[5][73] = -6'sd1;
    assign layer_1_weights[5][74] = 6'sd2;
    assign layer_1_weights[5][75] = 6'sd1;
    assign layer_1_weights[5][76] = 6'sd1;
    assign layer_1_weights[5][77] = -6'sd3;
    assign layer_1_weights[5][78] = -6'sd4;
    assign layer_1_weights[5][79] = 6'sd7;
    assign layer_1_weights[5][80] = 6'sd7;
    assign layer_1_weights[5][81] = 6'sd1;
    assign layer_1_weights[5][82] = 6'sd3;
    assign layer_1_weights[5][83] = 6'sd2;
    assign layer_1_weights[5][84] = -6'sd2;
    assign layer_1_weights[5][85] = 6'sd1;
    assign layer_1_weights[5][86] = 6'sd5;
    assign layer_1_weights[5][87] = 6'sd6;
    assign layer_1_weights[5][88] = 6'sd3;
    assign layer_1_weights[5][89] = -6'sd1;
    assign layer_1_weights[5][90] = 6'sd7;
    assign layer_1_weights[5][91] = 6'sd8;
    assign layer_1_weights[5][92] = 6'sd4;
    assign layer_1_weights[5][93] = 6'sd0;
    assign layer_1_weights[5][94] = 6'sd0;
    assign layer_1_weights[5][95] = -6'sd4;
    assign layer_1_weights[5][96] = 6'sd6;
    assign layer_1_weights[5][97] = 6'sd2;
    assign layer_1_weights[5][98] = -6'sd6;
    assign layer_1_weights[5][99] = -6'sd2;
    assign layer_1_weights[5][100] = 6'sd1;
    assign layer_1_weights[5][101] = 6'sd2;
    assign layer_1_weights[5][102] = 6'sd4;
    assign layer_1_weights[5][103] = 6'sd0;
    assign layer_1_weights[5][104] = -6'sd7;
    assign layer_1_weights[5][105] = -6'sd4;
    assign layer_1_weights[5][106] = -6'sd3;
    assign layer_1_weights[5][107] = 6'sd15;
    assign layer_1_weights[5][108] = -6'sd4;
    assign layer_1_weights[5][109] = 6'sd1;
    assign layer_1_weights[5][110] = -6'sd1;
    assign layer_1_weights[5][111] = -6'sd2;
    assign layer_1_weights[5][112] = -6'sd3;
    assign layer_1_weights[5][113] = -6'sd5;
    assign layer_1_weights[5][114] = -6'sd7;
    assign layer_1_weights[5][115] = -6'sd5;
    assign layer_1_weights[5][116] = -6'sd9;
    assign layer_1_weights[5][117] = -6'sd6;
    assign layer_1_weights[5][118] = -6'sd1;
    assign layer_1_weights[5][119] = -6'sd3;
    assign layer_1_weights[5][120] = -6'sd1;
    assign layer_1_weights[5][121] = 6'sd5;
    assign layer_1_weights[5][122] = 6'sd0;
    assign layer_1_weights[5][123] = -6'sd2;
    assign layer_1_weights[5][124] = -6'sd5;
    assign layer_1_weights[5][125] = -6'sd7;
    assign layer_1_weights[5][126] = -6'sd4;
    assign layer_1_weights[5][127] = -6'sd4;
    assign layer_1_weights[5][128] = -6'sd4;
    assign layer_1_weights[5][129] = -6'sd4;
    assign layer_1_weights[5][130] = -6'sd3;
    assign layer_1_weights[5][131] = 6'sd3;
    assign layer_1_weights[5][132] = -6'sd2;
    assign layer_1_weights[5][133] = 6'sd6;
    assign layer_1_weights[5][134] = 6'sd2;
    assign layer_1_weights[5][135] = 6'sd3;
    assign layer_1_weights[5][136] = -6'sd3;
    assign layer_1_weights[5][137] = 6'sd3;
    assign layer_1_weights[5][138] = 6'sd5;
    assign layer_1_weights[5][139] = 6'sd1;
    assign layer_1_weights[5][140] = -6'sd2;
    assign layer_1_weights[5][141] = 6'sd0;
    assign layer_1_weights[5][142] = 6'sd0;
    assign layer_1_weights[5][143] = 6'sd0;
    assign layer_1_biases[5] = 6'sd2;
    assign layer_1_weights[6][0] = 6'sd2;
    assign layer_1_weights[6][1] = 6'sd0;
    assign layer_1_weights[6][2] = -6'sd2;
    assign layer_1_weights[6][3] = -6'sd9;
    assign layer_1_weights[6][4] = -6'sd10;
    assign layer_1_weights[6][5] = -6'sd14;
    assign layer_1_weights[6][6] = -6'sd11;
    assign layer_1_weights[6][7] = -6'sd9;
    assign layer_1_weights[6][8] = -6'sd4;
    assign layer_1_weights[6][9] = -6'sd8;
    assign layer_1_weights[6][10] = -6'sd1;
    assign layer_1_weights[6][11] = -6'sd1;
    assign layer_1_weights[6][12] = -6'sd1;
    assign layer_1_weights[6][13] = 6'sd1;
    assign layer_1_weights[6][14] = 6'sd0;
    assign layer_1_weights[6][15] = -6'sd3;
    assign layer_1_weights[6][16] = -6'sd4;
    assign layer_1_weights[6][17] = -6'sd6;
    assign layer_1_weights[6][18] = -6'sd2;
    assign layer_1_weights[6][19] = -6'sd1;
    assign layer_1_weights[6][20] = 6'sd1;
    assign layer_1_weights[6][21] = 6'sd1;
    assign layer_1_weights[6][22] = 6'sd3;
    assign layer_1_weights[6][23] = 6'sd1;
    assign layer_1_weights[6][24] = -6'sd1;
    assign layer_1_weights[6][25] = -6'sd8;
    assign layer_1_weights[6][26] = 6'sd0;
    assign layer_1_weights[6][27] = 6'sd0;
    assign layer_1_weights[6][28] = 6'sd4;
    assign layer_1_weights[6][29] = 6'sd0;
    assign layer_1_weights[6][30] = 6'sd0;
    assign layer_1_weights[6][31] = -6'sd1;
    assign layer_1_weights[6][32] = -6'sd1;
    assign layer_1_weights[6][33] = 6'sd1;
    assign layer_1_weights[6][34] = -6'sd1;
    assign layer_1_weights[6][35] = 6'sd4;
    assign layer_1_weights[6][36] = -6'sd1;
    assign layer_1_weights[6][37] = 6'sd1;
    assign layer_1_weights[6][38] = -6'sd1;
    assign layer_1_weights[6][39] = 6'sd2;
    assign layer_1_weights[6][40] = 6'sd1;
    assign layer_1_weights[6][41] = 6'sd1;
    assign layer_1_weights[6][42] = -6'sd1;
    assign layer_1_weights[6][43] = -6'sd1;
    assign layer_1_weights[6][44] = 6'sd0;
    assign layer_1_weights[6][45] = -6'sd3;
    assign layer_1_weights[6][46] = 6'sd1;
    assign layer_1_weights[6][47] = 6'sd6;
    assign layer_1_weights[6][48] = -6'sd4;
    assign layer_1_weights[6][49] = -6'sd3;
    assign layer_1_weights[6][50] = 6'sd3;
    assign layer_1_weights[6][51] = 6'sd4;
    assign layer_1_weights[6][52] = 6'sd1;
    assign layer_1_weights[6][53] = -6'sd2;
    assign layer_1_weights[6][54] = -6'sd6;
    assign layer_1_weights[6][55] = -6'sd3;
    assign layer_1_weights[6][56] = 6'sd0;
    assign layer_1_weights[6][57] = 6'sd4;
    assign layer_1_weights[6][58] = 6'sd7;
    assign layer_1_weights[6][59] = 6'sd4;
    assign layer_1_weights[6][60] = -6'sd1;
    assign layer_1_weights[6][61] = -6'sd1;
    assign layer_1_weights[6][62] = 6'sd0;
    assign layer_1_weights[6][63] = 6'sd5;
    assign layer_1_weights[6][64] = 6'sd6;
    assign layer_1_weights[6][65] = 6'sd5;
    assign layer_1_weights[6][66] = -6'sd2;
    assign layer_1_weights[6][67] = 6'sd1;
    assign layer_1_weights[6][68] = -6'sd1;
    assign layer_1_weights[6][69] = 6'sd1;
    assign layer_1_weights[6][70] = 6'sd5;
    assign layer_1_weights[6][71] = -6'sd1;
    assign layer_1_weights[6][72] = -6'sd3;
    assign layer_1_weights[6][73] = -6'sd6;
    assign layer_1_weights[6][74] = 6'sd0;
    assign layer_1_weights[6][75] = 6'sd2;
    assign layer_1_weights[6][76] = 6'sd8;
    assign layer_1_weights[6][77] = 6'sd13;
    assign layer_1_weights[6][78] = 6'sd5;
    assign layer_1_weights[6][79] = -6'sd1;
    assign layer_1_weights[6][80] = -6'sd2;
    assign layer_1_weights[6][81] = -6'sd3;
    assign layer_1_weights[6][82] = 6'sd1;
    assign layer_1_weights[6][83] = -6'sd1;
    assign layer_1_weights[6][84] = -6'sd1;
    assign layer_1_weights[6][85] = -6'sd11;
    assign layer_1_weights[6][86] = -6'sd4;
    assign layer_1_weights[6][87] = -6'sd6;
    assign layer_1_weights[6][88] = -6'sd5;
    assign layer_1_weights[6][89] = -6'sd2;
    assign layer_1_weights[6][90] = 6'sd0;
    assign layer_1_weights[6][91] = -6'sd1;
    assign layer_1_weights[6][92] = -6'sd2;
    assign layer_1_weights[6][93] = -6'sd1;
    assign layer_1_weights[6][94] = 6'sd2;
    assign layer_1_weights[6][95] = -6'sd3;
    assign layer_1_weights[6][96] = 6'sd0;
    assign layer_1_weights[6][97] = -6'sd3;
    assign layer_1_weights[6][98] = -6'sd1;
    assign layer_1_weights[6][99] = -6'sd1;
    assign layer_1_weights[6][100] = -6'sd7;
    assign layer_1_weights[6][101] = -6'sd4;
    assign layer_1_weights[6][102] = -6'sd1;
    assign layer_1_weights[6][103] = 6'sd0;
    assign layer_1_weights[6][104] = -6'sd1;
    assign layer_1_weights[6][105] = 6'sd1;
    assign layer_1_weights[6][106] = 6'sd0;
    assign layer_1_weights[6][107] = -6'sd11;
    assign layer_1_weights[6][108] = 6'sd0;
    assign layer_1_weights[6][109] = 6'sd3;
    assign layer_1_weights[6][110] = 6'sd0;
    assign layer_1_weights[6][111] = 6'sd4;
    assign layer_1_weights[6][112] = 6'sd2;
    assign layer_1_weights[6][113] = 6'sd1;
    assign layer_1_weights[6][114] = -6'sd2;
    assign layer_1_weights[6][115] = -6'sd3;
    assign layer_1_weights[6][116] = 6'sd0;
    assign layer_1_weights[6][117] = 6'sd0;
    assign layer_1_weights[6][118] = 6'sd0;
    assign layer_1_weights[6][119] = 6'sd4;
    assign layer_1_weights[6][120] = 6'sd1;
    assign layer_1_weights[6][121] = 6'sd4;
    assign layer_1_weights[6][122] = -6'sd1;
    assign layer_1_weights[6][123] = 6'sd2;
    assign layer_1_weights[6][124] = 6'sd3;
    assign layer_1_weights[6][125] = 6'sd2;
    assign layer_1_weights[6][126] = 6'sd0;
    assign layer_1_weights[6][127] = -6'sd1;
    assign layer_1_weights[6][128] = -6'sd1;
    assign layer_1_weights[6][129] = 6'sd0;
    assign layer_1_weights[6][130] = 6'sd1;
    assign layer_1_weights[6][131] = -6'sd5;
    assign layer_1_weights[6][132] = -6'sd1;
    assign layer_1_weights[6][133] = 6'sd1;
    assign layer_1_weights[6][134] = -6'sd6;
    assign layer_1_weights[6][135] = -6'sd2;
    assign layer_1_weights[6][136] = 6'sd1;
    assign layer_1_weights[6][137] = 6'sd0;
    assign layer_1_weights[6][138] = 6'sd5;
    assign layer_1_weights[6][139] = 6'sd8;
    assign layer_1_weights[6][140] = 6'sd0;
    assign layer_1_weights[6][141] = 6'sd6;
    assign layer_1_weights[6][142] = 6'sd1;
    assign layer_1_weights[6][143] = 6'sd0;
    assign layer_1_biases[6] = -6'sd1;
    assign layer_1_weights[7][0] = -6'sd2;
    assign layer_1_weights[7][1] = 6'sd1;
    assign layer_1_weights[7][2] = 6'sd3;
    assign layer_1_weights[7][3] = 6'sd13;
    assign layer_1_weights[7][4] = 6'sd16;
    assign layer_1_weights[7][5] = 6'sd4;
    assign layer_1_weights[7][6] = -6'sd3;
    assign layer_1_weights[7][7] = 6'sd5;
    assign layer_1_weights[7][8] = -6'sd2;
    assign layer_1_weights[7][9] = 6'sd11;
    assign layer_1_weights[7][10] = 6'sd1;
    assign layer_1_weights[7][11] = 6'sd1;
    assign layer_1_weights[7][12] = 6'sd0;
    assign layer_1_weights[7][13] = 6'sd2;
    assign layer_1_weights[7][14] = 6'sd7;
    assign layer_1_weights[7][15] = 6'sd1;
    assign layer_1_weights[7][16] = 6'sd0;
    assign layer_1_weights[7][17] = 6'sd1;
    assign layer_1_weights[7][18] = -6'sd2;
    assign layer_1_weights[7][19] = -6'sd1;
    assign layer_1_weights[7][20] = -6'sd2;
    assign layer_1_weights[7][21] = 6'sd1;
    assign layer_1_weights[7][22] = 6'sd0;
    assign layer_1_weights[7][23] = -6'sd3;
    assign layer_1_weights[7][24] = 6'sd0;
    assign layer_1_weights[7][25] = 6'sd1;
    assign layer_1_weights[7][26] = 6'sd4;
    assign layer_1_weights[7][27] = -6'sd2;
    assign layer_1_weights[7][28] = 6'sd0;
    assign layer_1_weights[7][29] = -6'sd1;
    assign layer_1_weights[7][30] = -6'sd1;
    assign layer_1_weights[7][31] = -6'sd3;
    assign layer_1_weights[7][32] = -6'sd2;
    assign layer_1_weights[7][33] = 6'sd0;
    assign layer_1_weights[7][34] = 6'sd0;
    assign layer_1_weights[7][35] = 6'sd2;
    assign layer_1_weights[7][36] = 6'sd4;
    assign layer_1_weights[7][37] = -6'sd4;
    assign layer_1_weights[7][38] = -6'sd4;
    assign layer_1_weights[7][39] = -6'sd4;
    assign layer_1_weights[7][40] = -6'sd4;
    assign layer_1_weights[7][41] = -6'sd2;
    assign layer_1_weights[7][42] = -6'sd2;
    assign layer_1_weights[7][43] = -6'sd4;
    assign layer_1_weights[7][44] = 6'sd0;
    assign layer_1_weights[7][45] = 6'sd1;
    assign layer_1_weights[7][46] = 6'sd2;
    assign layer_1_weights[7][47] = 6'sd5;
    assign layer_1_weights[7][48] = -6'sd1;
    assign layer_1_weights[7][49] = -6'sd9;
    assign layer_1_weights[7][50] = -6'sd6;
    assign layer_1_weights[7][51] = -6'sd7;
    assign layer_1_weights[7][52] = -6'sd6;
    assign layer_1_weights[7][53] = -6'sd1;
    assign layer_1_weights[7][54] = -6'sd1;
    assign layer_1_weights[7][55] = -6'sd4;
    assign layer_1_weights[7][56] = -6'sd2;
    assign layer_1_weights[7][57] = 6'sd0;
    assign layer_1_weights[7][58] = -6'sd3;
    assign layer_1_weights[7][59] = -6'sd6;
    assign layer_1_weights[7][60] = 6'sd0;
    assign layer_1_weights[7][61] = -6'sd4;
    assign layer_1_weights[7][62] = -6'sd3;
    assign layer_1_weights[7][63] = 6'sd0;
    assign layer_1_weights[7][64] = 6'sd5;
    assign layer_1_weights[7][65] = 6'sd9;
    assign layer_1_weights[7][66] = -6'sd1;
    assign layer_1_weights[7][67] = -6'sd2;
    assign layer_1_weights[7][68] = -6'sd2;
    assign layer_1_weights[7][69] = -6'sd2;
    assign layer_1_weights[7][70] = 6'sd0;
    assign layer_1_weights[7][71] = 6'sd1;
    assign layer_1_weights[7][72] = 6'sd2;
    assign layer_1_weights[7][73] = 6'sd2;
    assign layer_1_weights[7][74] = 6'sd4;
    assign layer_1_weights[7][75] = 6'sd6;
    assign layer_1_weights[7][76] = 6'sd6;
    assign layer_1_weights[7][77] = 6'sd6;
    assign layer_1_weights[7][78] = 6'sd5;
    assign layer_1_weights[7][79] = 6'sd1;
    assign layer_1_weights[7][80] = 6'sd1;
    assign layer_1_weights[7][81] = 6'sd1;
    assign layer_1_weights[7][82] = 6'sd2;
    assign layer_1_weights[7][83] = 6'sd8;
    assign layer_1_weights[7][84] = 6'sd1;
    assign layer_1_weights[7][85] = 6'sd7;
    assign layer_1_weights[7][86] = 6'sd3;
    assign layer_1_weights[7][87] = 6'sd3;
    assign layer_1_weights[7][88] = 6'sd0;
    assign layer_1_weights[7][89] = 6'sd0;
    assign layer_1_weights[7][90] = 6'sd4;
    assign layer_1_weights[7][91] = 6'sd5;
    assign layer_1_weights[7][92] = 6'sd6;
    assign layer_1_weights[7][93] = 6'sd7;
    assign layer_1_weights[7][94] = 6'sd5;
    assign layer_1_weights[7][95] = 6'sd9;
    assign layer_1_weights[7][96] = 6'sd0;
    assign layer_1_weights[7][97] = -6'sd1;
    assign layer_1_weights[7][98] = -6'sd3;
    assign layer_1_weights[7][99] = 6'sd1;
    assign layer_1_weights[7][100] = -6'sd1;
    assign layer_1_weights[7][101] = -6'sd2;
    assign layer_1_weights[7][102] = 6'sd5;
    assign layer_1_weights[7][103] = 6'sd3;
    assign layer_1_weights[7][104] = 6'sd3;
    assign layer_1_weights[7][105] = 6'sd1;
    assign layer_1_weights[7][106] = -6'sd1;
    assign layer_1_weights[7][107] = 6'sd7;
    assign layer_1_weights[7][108] = -6'sd1;
    assign layer_1_weights[7][109] = -6'sd4;
    assign layer_1_weights[7][110] = -6'sd4;
    assign layer_1_weights[7][111] = -6'sd1;
    assign layer_1_weights[7][112] = -6'sd2;
    assign layer_1_weights[7][113] = -6'sd3;
    assign layer_1_weights[7][114] = -6'sd5;
    assign layer_1_weights[7][115] = -6'sd2;
    assign layer_1_weights[7][116] = -6'sd2;
    assign layer_1_weights[7][117] = -6'sd4;
    assign layer_1_weights[7][118] = -6'sd1;
    assign layer_1_weights[7][119] = -6'sd2;
    assign layer_1_weights[7][120] = 6'sd1;
    assign layer_1_weights[7][121] = 6'sd0;
    assign layer_1_weights[7][122] = 6'sd2;
    assign layer_1_weights[7][123] = -6'sd2;
    assign layer_1_weights[7][124] = 6'sd0;
    assign layer_1_weights[7][125] = 6'sd1;
    assign layer_1_weights[7][126] = 6'sd0;
    assign layer_1_weights[7][127] = -6'sd3;
    assign layer_1_weights[7][128] = -6'sd1;
    assign layer_1_weights[7][129] = 6'sd4;
    assign layer_1_weights[7][130] = -6'sd10;
    assign layer_1_weights[7][131] = 6'sd4;
    assign layer_1_weights[7][132] = -6'sd1;
    assign layer_1_weights[7][133] = -6'sd4;
    assign layer_1_weights[7][134] = -6'sd14;
    assign layer_1_weights[7][135] = -6'sd17;
    assign layer_1_weights[7][136] = -6'sd14;
    assign layer_1_weights[7][137] = -6'sd8;
    assign layer_1_weights[7][138] = -6'sd6;
    assign layer_1_weights[7][139] = -6'sd9;
    assign layer_1_weights[7][140] = -6'sd13;
    assign layer_1_weights[7][141] = -6'sd2;
    assign layer_1_weights[7][142] = 6'sd1;
    assign layer_1_weights[7][143] = -6'sd1;
    assign layer_1_biases[7] = 6'sd6;
    assign layer_1_weights[8][0] = -6'sd1;
    assign layer_1_weights[8][1] = 6'sd0;
    assign layer_1_weights[8][2] = 6'sd5;
    assign layer_1_weights[8][3] = 6'sd7;
    assign layer_1_weights[8][4] = 6'sd5;
    assign layer_1_weights[8][5] = 6'sd1;
    assign layer_1_weights[8][6] = 6'sd6;
    assign layer_1_weights[8][7] = 6'sd0;
    assign layer_1_weights[8][8] = 6'sd0;
    assign layer_1_weights[8][9] = 6'sd10;
    assign layer_1_weights[8][10] = 6'sd0;
    assign layer_1_weights[8][11] = -6'sd1;
    assign layer_1_weights[8][12] = -6'sd1;
    assign layer_1_weights[8][13] = 6'sd2;
    assign layer_1_weights[8][14] = 6'sd1;
    assign layer_1_weights[8][15] = 6'sd4;
    assign layer_1_weights[8][16] = 6'sd6;
    assign layer_1_weights[8][17] = 6'sd5;
    assign layer_1_weights[8][18] = 6'sd6;
    assign layer_1_weights[8][19] = 6'sd6;
    assign layer_1_weights[8][20] = 6'sd3;
    assign layer_1_weights[8][21] = 6'sd1;
    assign layer_1_weights[8][22] = -6'sd4;
    assign layer_1_weights[8][23] = 6'sd1;
    assign layer_1_weights[8][24] = 6'sd1;
    assign layer_1_weights[8][25] = -6'sd6;
    assign layer_1_weights[8][26] = 6'sd4;
    assign layer_1_weights[8][27] = 6'sd2;
    assign layer_1_weights[8][28] = 6'sd3;
    assign layer_1_weights[8][29] = 6'sd1;
    assign layer_1_weights[8][30] = 6'sd0;
    assign layer_1_weights[8][31] = -6'sd1;
    assign layer_1_weights[8][32] = -6'sd1;
    assign layer_1_weights[8][33] = 6'sd4;
    assign layer_1_weights[8][34] = 6'sd3;
    assign layer_1_weights[8][35] = 6'sd5;
    assign layer_1_weights[8][36] = -6'sd5;
    assign layer_1_weights[8][37] = 6'sd3;
    assign layer_1_weights[8][38] = -6'sd1;
    assign layer_1_weights[8][39] = 6'sd2;
    assign layer_1_weights[8][40] = 6'sd1;
    assign layer_1_weights[8][41] = -6'sd3;
    assign layer_1_weights[8][42] = -6'sd2;
    assign layer_1_weights[8][43] = 6'sd1;
    assign layer_1_weights[8][44] = 6'sd2;
    assign layer_1_weights[8][45] = 6'sd0;
    assign layer_1_weights[8][46] = 6'sd0;
    assign layer_1_weights[8][47] = 6'sd4;
    assign layer_1_weights[8][48] = -6'sd1;
    assign layer_1_weights[8][49] = 6'sd3;
    assign layer_1_weights[8][50] = -6'sd1;
    assign layer_1_weights[8][51] = -6'sd2;
    assign layer_1_weights[8][52] = 6'sd1;
    assign layer_1_weights[8][53] = 6'sd0;
    assign layer_1_weights[8][54] = 6'sd2;
    assign layer_1_weights[8][55] = -6'sd3;
    assign layer_1_weights[8][56] = -6'sd1;
    assign layer_1_weights[8][57] = 6'sd0;
    assign layer_1_weights[8][58] = 6'sd4;
    assign layer_1_weights[8][59] = 6'sd3;
    assign layer_1_weights[8][60] = -6'sd5;
    assign layer_1_weights[8][61] = -6'sd7;
    assign layer_1_weights[8][62] = 6'sd1;
    assign layer_1_weights[8][63] = 6'sd1;
    assign layer_1_weights[8][64] = 6'sd5;
    assign layer_1_weights[8][65] = 6'sd5;
    assign layer_1_weights[8][66] = 6'sd3;
    assign layer_1_weights[8][67] = 6'sd1;
    assign layer_1_weights[8][68] = 6'sd3;
    assign layer_1_weights[8][69] = 6'sd2;
    assign layer_1_weights[8][70] = -6'sd3;
    assign layer_1_weights[8][71] = -6'sd4;
    assign layer_1_weights[8][72] = 6'sd2;
    assign layer_1_weights[8][73] = 6'sd3;
    assign layer_1_weights[8][74] = 6'sd5;
    assign layer_1_weights[8][75] = 6'sd4;
    assign layer_1_weights[8][76] = 6'sd3;
    assign layer_1_weights[8][77] = 6'sd5;
    assign layer_1_weights[8][78] = 6'sd0;
    assign layer_1_weights[8][79] = -6'sd1;
    assign layer_1_weights[8][80] = -6'sd3;
    assign layer_1_weights[8][81] = -6'sd1;
    assign layer_1_weights[8][82] = 6'sd0;
    assign layer_1_weights[8][83] = -6'sd7;
    assign layer_1_weights[8][84] = 6'sd3;
    assign layer_1_weights[8][85] = 6'sd0;
    assign layer_1_weights[8][86] = 6'sd1;
    assign layer_1_weights[8][87] = -6'sd2;
    assign layer_1_weights[8][88] = 6'sd2;
    assign layer_1_weights[8][89] = 6'sd4;
    assign layer_1_weights[8][90] = 6'sd1;
    assign layer_1_weights[8][91] = 6'sd2;
    assign layer_1_weights[8][92] = -6'sd1;
    assign layer_1_weights[8][93] = 6'sd2;
    assign layer_1_weights[8][94] = 6'sd2;
    assign layer_1_weights[8][95] = -6'sd3;
    assign layer_1_weights[8][96] = 6'sd4;
    assign layer_1_weights[8][97] = -6'sd1;
    assign layer_1_weights[8][98] = -6'sd2;
    assign layer_1_weights[8][99] = 6'sd0;
    assign layer_1_weights[8][100] = 6'sd2;
    assign layer_1_weights[8][101] = 6'sd2;
    assign layer_1_weights[8][102] = 6'sd0;
    assign layer_1_weights[8][103] = 6'sd2;
    assign layer_1_weights[8][104] = 6'sd5;
    assign layer_1_weights[8][105] = 6'sd0;
    assign layer_1_weights[8][106] = -6'sd3;
    assign layer_1_weights[8][107] = -6'sd7;
    assign layer_1_weights[8][108] = -6'sd4;
    assign layer_1_weights[8][109] = 6'sd1;
    assign layer_1_weights[8][110] = 6'sd2;
    assign layer_1_weights[8][111] = -6'sd1;
    assign layer_1_weights[8][112] = -6'sd1;
    assign layer_1_weights[8][113] = 6'sd3;
    assign layer_1_weights[8][114] = 6'sd5;
    assign layer_1_weights[8][115] = 6'sd7;
    assign layer_1_weights[8][116] = 6'sd5;
    assign layer_1_weights[8][117] = -6'sd1;
    assign layer_1_weights[8][118] = -6'sd3;
    assign layer_1_weights[8][119] = 6'sd4;
    assign layer_1_weights[8][120] = -6'sd1;
    assign layer_1_weights[8][121] = -6'sd3;
    assign layer_1_weights[8][122] = -6'sd2;
    assign layer_1_weights[8][123] = 6'sd0;
    assign layer_1_weights[8][124] = 6'sd0;
    assign layer_1_weights[8][125] = 6'sd6;
    assign layer_1_weights[8][126] = 6'sd6;
    assign layer_1_weights[8][127] = 6'sd8;
    assign layer_1_weights[8][128] = 6'sd0;
    assign layer_1_weights[8][129] = -6'sd3;
    assign layer_1_weights[8][130] = -6'sd7;
    assign layer_1_weights[8][131] = -6'sd5;
    assign layer_1_weights[8][132] = 6'sd2;
    assign layer_1_weights[8][133] = -6'sd3;
    assign layer_1_weights[8][134] = 6'sd0;
    assign layer_1_weights[8][135] = -6'sd3;
    assign layer_1_weights[8][136] = 6'sd0;
    assign layer_1_weights[8][137] = -6'sd2;
    assign layer_1_weights[8][138] = -6'sd6;
    assign layer_1_weights[8][139] = -6'sd5;
    assign layer_1_weights[8][140] = 6'sd0;
    assign layer_1_weights[8][141] = -6'sd2;
    assign layer_1_weights[8][142] = 6'sd0;
    assign layer_1_weights[8][143] = -6'sd2;
    assign layer_1_biases[8] = -6'sd4;
    assign layer_1_weights[9][0] = -6'sd1;
    assign layer_1_weights[9][1] = 6'sd1;
    assign layer_1_weights[9][2] = 6'sd0;
    assign layer_1_weights[9][3] = 6'sd0;
    assign layer_1_weights[9][4] = -6'sd1;
    assign layer_1_weights[9][5] = 6'sd1;
    assign layer_1_weights[9][6] = 6'sd3;
    assign layer_1_weights[9][7] = -6'sd7;
    assign layer_1_weights[9][8] = 6'sd5;
    assign layer_1_weights[9][9] = -6'sd1;
    assign layer_1_weights[9][10] = -6'sd1;
    assign layer_1_weights[9][11] = 6'sd1;
    assign layer_1_weights[9][12] = -6'sd2;
    assign layer_1_weights[9][13] = 6'sd0;
    assign layer_1_weights[9][14] = -6'sd8;
    assign layer_1_weights[9][15] = -6'sd6;
    assign layer_1_weights[9][16] = -6'sd7;
    assign layer_1_weights[9][17] = -6'sd3;
    assign layer_1_weights[9][18] = -6'sd3;
    assign layer_1_weights[9][19] = 6'sd0;
    assign layer_1_weights[9][20] = 6'sd3;
    assign layer_1_weights[9][21] = 6'sd0;
    assign layer_1_weights[9][22] = -6'sd11;
    assign layer_1_weights[9][23] = -6'sd1;
    assign layer_1_weights[9][24] = 6'sd1;
    assign layer_1_weights[9][25] = -6'sd5;
    assign layer_1_weights[9][26] = -6'sd3;
    assign layer_1_weights[9][27] = -6'sd1;
    assign layer_1_weights[9][28] = 6'sd0;
    assign layer_1_weights[9][29] = 6'sd2;
    assign layer_1_weights[9][30] = 6'sd0;
    assign layer_1_weights[9][31] = -6'sd4;
    assign layer_1_weights[9][32] = 6'sd1;
    assign layer_1_weights[9][33] = 6'sd1;
    assign layer_1_weights[9][34] = -6'sd1;
    assign layer_1_weights[9][35] = -6'sd3;
    assign layer_1_weights[9][36] = 6'sd4;
    assign layer_1_weights[9][37] = 6'sd3;
    assign layer_1_weights[9][38] = -6'sd2;
    assign layer_1_weights[9][39] = -6'sd2;
    assign layer_1_weights[9][40] = -6'sd2;
    assign layer_1_weights[9][41] = 6'sd5;
    assign layer_1_weights[9][42] = 6'sd2;
    assign layer_1_weights[9][43] = 6'sd1;
    assign layer_1_weights[9][44] = 6'sd0;
    assign layer_1_weights[9][45] = 6'sd1;
    assign layer_1_weights[9][46] = 6'sd2;
    assign layer_1_weights[9][47] = -6'sd3;
    assign layer_1_weights[9][48] = 6'sd11;
    assign layer_1_weights[9][49] = 6'sd6;
    assign layer_1_weights[9][50] = 6'sd3;
    assign layer_1_weights[9][51] = 6'sd2;
    assign layer_1_weights[9][52] = 6'sd5;
    assign layer_1_weights[9][53] = 6'sd6;
    assign layer_1_weights[9][54] = 6'sd4;
    assign layer_1_weights[9][55] = 6'sd2;
    assign layer_1_weights[9][56] = 6'sd3;
    assign layer_1_weights[9][57] = 6'sd0;
    assign layer_1_weights[9][58] = 6'sd1;
    assign layer_1_weights[9][59] = 6'sd4;
    assign layer_1_weights[9][60] = 6'sd13;
    assign layer_1_weights[9][61] = -6'sd3;
    assign layer_1_weights[9][62] = 6'sd3;
    assign layer_1_weights[9][63] = 6'sd2;
    assign layer_1_weights[9][64] = 6'sd3;
    assign layer_1_weights[9][65] = -6'sd4;
    assign layer_1_weights[9][66] = -6'sd9;
    assign layer_1_weights[9][67] = -6'sd4;
    assign layer_1_weights[9][68] = 6'sd0;
    assign layer_1_weights[9][69] = -6'sd2;
    assign layer_1_weights[9][70] = -6'sd1;
    assign layer_1_weights[9][71] = 6'sd4;
    assign layer_1_weights[9][72] = 6'sd1;
    assign layer_1_weights[9][73] = -6'sd4;
    assign layer_1_weights[9][74] = -6'sd2;
    assign layer_1_weights[9][75] = -6'sd1;
    assign layer_1_weights[9][76] = -6'sd3;
    assign layer_1_weights[9][77] = -6'sd10;
    assign layer_1_weights[9][78] = -6'sd6;
    assign layer_1_weights[9][79] = 6'sd0;
    assign layer_1_weights[9][80] = -6'sd6;
    assign layer_1_weights[9][81] = -6'sd3;
    assign layer_1_weights[9][82] = -6'sd2;
    assign layer_1_weights[9][83] = 6'sd6;
    assign layer_1_weights[9][84] = -6'sd3;
    assign layer_1_weights[9][85] = -6'sd1;
    assign layer_1_weights[9][86] = -6'sd2;
    assign layer_1_weights[9][87] = -6'sd3;
    assign layer_1_weights[9][88] = -6'sd6;
    assign layer_1_weights[9][89] = -6'sd6;
    assign layer_1_weights[9][90] = -6'sd1;
    assign layer_1_weights[9][91] = -6'sd1;
    assign layer_1_weights[9][92] = -6'sd3;
    assign layer_1_weights[9][93] = -6'sd1;
    assign layer_1_weights[9][94] = -6'sd2;
    assign layer_1_weights[9][95] = 6'sd16;
    assign layer_1_weights[9][96] = -6'sd4;
    assign layer_1_weights[9][97] = 6'sd0;
    assign layer_1_weights[9][98] = 6'sd3;
    assign layer_1_weights[9][99] = -6'sd1;
    assign layer_1_weights[9][100] = 6'sd0;
    assign layer_1_weights[9][101] = 6'sd1;
    assign layer_1_weights[9][102] = 6'sd4;
    assign layer_1_weights[9][103] = 6'sd2;
    assign layer_1_weights[9][104] = 6'sd4;
    assign layer_1_weights[9][105] = 6'sd3;
    assign layer_1_weights[9][106] = 6'sd3;
    assign layer_1_weights[9][107] = 6'sd7;
    assign layer_1_weights[9][108] = -6'sd2;
    assign layer_1_weights[9][109] = 6'sd1;
    assign layer_1_weights[9][110] = 6'sd5;
    assign layer_1_weights[9][111] = 6'sd5;
    assign layer_1_weights[9][112] = 6'sd5;
    assign layer_1_weights[9][113] = 6'sd2;
    assign layer_1_weights[9][114] = 6'sd4;
    assign layer_1_weights[9][115] = 6'sd5;
    assign layer_1_weights[9][116] = 6'sd3;
    assign layer_1_weights[9][117] = 6'sd1;
    assign layer_1_weights[9][118] = 6'sd10;
    assign layer_1_weights[9][119] = 6'sd6;
    assign layer_1_weights[9][120] = -6'sd1;
    assign layer_1_weights[9][121] = 6'sd1;
    assign layer_1_weights[9][122] = 6'sd3;
    assign layer_1_weights[9][123] = 6'sd2;
    assign layer_1_weights[9][124] = 6'sd0;
    assign layer_1_weights[9][125] = 6'sd1;
    assign layer_1_weights[9][126] = 6'sd0;
    assign layer_1_weights[9][127] = -6'sd1;
    assign layer_1_weights[9][128] = 6'sd0;
    assign layer_1_weights[9][129] = 6'sd0;
    assign layer_1_weights[9][130] = 6'sd2;
    assign layer_1_weights[9][131] = 6'sd1;
    assign layer_1_weights[9][132] = 6'sd0;
    assign layer_1_weights[9][133] = 6'sd0;
    assign layer_1_weights[9][134] = 6'sd1;
    assign layer_1_weights[9][135] = 6'sd2;
    assign layer_1_weights[9][136] = -6'sd1;
    assign layer_1_weights[9][137] = -6'sd2;
    assign layer_1_weights[9][138] = 6'sd2;
    assign layer_1_weights[9][139] = -6'sd2;
    assign layer_1_weights[9][140] = -6'sd2;
    assign layer_1_weights[9][141] = 6'sd0;
    assign layer_1_weights[9][142] = 6'sd1;
    assign layer_1_weights[9][143] = 6'sd1;
    assign layer_1_biases[9] = 6'sd2;
    assign layer_1_weights[10][0] = 6'sd0;
    assign layer_1_weights[10][1] = 6'sd2;
    assign layer_1_weights[10][2] = 6'sd4;
    assign layer_1_weights[10][3] = 6'sd7;
    assign layer_1_weights[10][4] = 6'sd3;
    assign layer_1_weights[10][5] = 6'sd1;
    assign layer_1_weights[10][6] = 6'sd2;
    assign layer_1_weights[10][7] = 6'sd7;
    assign layer_1_weights[10][8] = -6'sd2;
    assign layer_1_weights[10][9] = 6'sd9;
    assign layer_1_weights[10][10] = 6'sd2;
    assign layer_1_weights[10][11] = -6'sd1;
    assign layer_1_weights[10][12] = 6'sd1;
    assign layer_1_weights[10][13] = 6'sd0;
    assign layer_1_weights[10][14] = 6'sd1;
    assign layer_1_weights[10][15] = 6'sd1;
    assign layer_1_weights[10][16] = 6'sd3;
    assign layer_1_weights[10][17] = 6'sd2;
    assign layer_1_weights[10][18] = -6'sd2;
    assign layer_1_weights[10][19] = 6'sd0;
    assign layer_1_weights[10][20] = -6'sd3;
    assign layer_1_weights[10][21] = 6'sd5;
    assign layer_1_weights[10][22] = -6'sd11;
    assign layer_1_weights[10][23] = -6'sd2;
    assign layer_1_weights[10][24] = 6'sd0;
    assign layer_1_weights[10][25] = -6'sd2;
    assign layer_1_weights[10][26] = -6'sd2;
    assign layer_1_weights[10][27] = 6'sd0;
    assign layer_1_weights[10][28] = 6'sd0;
    assign layer_1_weights[10][29] = 6'sd2;
    assign layer_1_weights[10][30] = 6'sd0;
    assign layer_1_weights[10][31] = 6'sd2;
    assign layer_1_weights[10][32] = 6'sd1;
    assign layer_1_weights[10][33] = -6'sd1;
    assign layer_1_weights[10][34] = -6'sd5;
    assign layer_1_weights[10][35] = 6'sd0;
    assign layer_1_weights[10][36] = 6'sd0;
    assign layer_1_weights[10][37] = 6'sd1;
    assign layer_1_weights[10][38] = 6'sd0;
    assign layer_1_weights[10][39] = 6'sd0;
    assign layer_1_weights[10][40] = 6'sd6;
    assign layer_1_weights[10][41] = 6'sd3;
    assign layer_1_weights[10][42] = -6'sd1;
    assign layer_1_weights[10][43] = -6'sd3;
    assign layer_1_weights[10][44] = -6'sd1;
    assign layer_1_weights[10][45] = 6'sd3;
    assign layer_1_weights[10][46] = -6'sd1;
    assign layer_1_weights[10][47] = -6'sd9;
    assign layer_1_weights[10][48] = 6'sd4;
    assign layer_1_weights[10][49] = -6'sd3;
    assign layer_1_weights[10][50] = -6'sd2;
    assign layer_1_weights[10][51] = 6'sd1;
    assign layer_1_weights[10][52] = 6'sd5;
    assign layer_1_weights[10][53] = -6'sd6;
    assign layer_1_weights[10][54] = -6'sd2;
    assign layer_1_weights[10][55] = 6'sd0;
    assign layer_1_weights[10][56] = -6'sd1;
    assign layer_1_weights[10][57] = -6'sd1;
    assign layer_1_weights[10][58] = -6'sd3;
    assign layer_1_weights[10][59] = -6'sd4;
    assign layer_1_weights[10][60] = 6'sd2;
    assign layer_1_weights[10][61] = 6'sd1;
    assign layer_1_weights[10][62] = 6'sd3;
    assign layer_1_weights[10][63] = 6'sd5;
    assign layer_1_weights[10][64] = 6'sd0;
    assign layer_1_weights[10][65] = -6'sd7;
    assign layer_1_weights[10][66] = -6'sd3;
    assign layer_1_weights[10][67] = 6'sd5;
    assign layer_1_weights[10][68] = 6'sd0;
    assign layer_1_weights[10][69] = 6'sd4;
    assign layer_1_weights[10][70] = 6'sd4;
    assign layer_1_weights[10][71] = 6'sd0;
    assign layer_1_weights[10][72] = 6'sd1;
    assign layer_1_weights[10][73] = 6'sd6;
    assign layer_1_weights[10][74] = 6'sd5;
    assign layer_1_weights[10][75] = 6'sd5;
    assign layer_1_weights[10][76] = -6'sd1;
    assign layer_1_weights[10][77] = -6'sd6;
    assign layer_1_weights[10][78] = 6'sd0;
    assign layer_1_weights[10][79] = -6'sd4;
    assign layer_1_weights[10][80] = 6'sd1;
    assign layer_1_weights[10][81] = 6'sd5;
    assign layer_1_weights[10][82] = 6'sd7;
    assign layer_1_weights[10][83] = -6'sd4;
    assign layer_1_weights[10][84] = -6'sd2;
    assign layer_1_weights[10][85] = -6'sd1;
    assign layer_1_weights[10][86] = 6'sd2;
    assign layer_1_weights[10][87] = 6'sd4;
    assign layer_1_weights[10][88] = 6'sd2;
    assign layer_1_weights[10][89] = -6'sd4;
    assign layer_1_weights[10][90] = -6'sd7;
    assign layer_1_weights[10][91] = -6'sd1;
    assign layer_1_weights[10][92] = 6'sd4;
    assign layer_1_weights[10][93] = 6'sd0;
    assign layer_1_weights[10][94] = 6'sd0;
    assign layer_1_weights[10][95] = -6'sd1;
    assign layer_1_weights[10][96] = -6'sd5;
    assign layer_1_weights[10][97] = -6'sd1;
    assign layer_1_weights[10][98] = -6'sd2;
    assign layer_1_weights[10][99] = 6'sd1;
    assign layer_1_weights[10][100] = 6'sd2;
    assign layer_1_weights[10][101] = -6'sd1;
    assign layer_1_weights[10][102] = -6'sd1;
    assign layer_1_weights[10][103] = 6'sd8;
    assign layer_1_weights[10][104] = 6'sd3;
    assign layer_1_weights[10][105] = 6'sd0;
    assign layer_1_weights[10][106] = -6'sd2;
    assign layer_1_weights[10][107] = -6'sd11;
    assign layer_1_weights[10][108] = -6'sd6;
    assign layer_1_weights[10][109] = -6'sd4;
    assign layer_1_weights[10][110] = -6'sd4;
    assign layer_1_weights[10][111] = -6'sd3;
    assign layer_1_weights[10][112] = -6'sd4;
    assign layer_1_weights[10][113] = -6'sd1;
    assign layer_1_weights[10][114] = 6'sd6;
    assign layer_1_weights[10][115] = 6'sd5;
    assign layer_1_weights[10][116] = 6'sd2;
    assign layer_1_weights[10][117] = -6'sd2;
    assign layer_1_weights[10][118] = 6'sd1;
    assign layer_1_weights[10][119] = 6'sd4;
    assign layer_1_weights[10][120] = -6'sd1;
    assign layer_1_weights[10][121] = 6'sd3;
    assign layer_1_weights[10][122] = -6'sd3;
    assign layer_1_weights[10][123] = -6'sd4;
    assign layer_1_weights[10][124] = -6'sd2;
    assign layer_1_weights[10][125] = 6'sd0;
    assign layer_1_weights[10][126] = 6'sd7;
    assign layer_1_weights[10][127] = 6'sd6;
    assign layer_1_weights[10][128] = 6'sd3;
    assign layer_1_weights[10][129] = -6'sd2;
    assign layer_1_weights[10][130] = -6'sd5;
    assign layer_1_weights[10][131] = -6'sd4;
    assign layer_1_weights[10][132] = -6'sd1;
    assign layer_1_weights[10][133] = 6'sd1;
    assign layer_1_weights[10][134] = -6'sd5;
    assign layer_1_weights[10][135] = -6'sd5;
    assign layer_1_weights[10][136] = 6'sd4;
    assign layer_1_weights[10][137] = 6'sd0;
    assign layer_1_weights[10][138] = 6'sd5;
    assign layer_1_weights[10][139] = -6'sd1;
    assign layer_1_weights[10][140] = 6'sd4;
    assign layer_1_weights[10][141] = 6'sd7;
    assign layer_1_weights[10][142] = -6'sd1;
    assign layer_1_weights[10][143] = -6'sd1;
    assign layer_1_biases[10] = -6'sd4;
    assign layer_1_weights[11][0] = 6'sd1;
    assign layer_1_weights[11][1] = -6'sd2;
    assign layer_1_weights[11][2] = 6'sd0;
    assign layer_1_weights[11][3] = 6'sd5;
    assign layer_1_weights[11][4] = 6'sd4;
    assign layer_1_weights[11][5] = 6'sd5;
    assign layer_1_weights[11][6] = 6'sd6;
    assign layer_1_weights[11][7] = 6'sd2;
    assign layer_1_weights[11][8] = 6'sd2;
    assign layer_1_weights[11][9] = 6'sd7;
    assign layer_1_weights[11][10] = -6'sd2;
    assign layer_1_weights[11][11] = -6'sd1;
    assign layer_1_weights[11][12] = 6'sd1;
    assign layer_1_weights[11][13] = 6'sd0;
    assign layer_1_weights[11][14] = -6'sd4;
    assign layer_1_weights[11][15] = 6'sd2;
    assign layer_1_weights[11][16] = 6'sd3;
    assign layer_1_weights[11][17] = 6'sd5;
    assign layer_1_weights[11][18] = 6'sd7;
    assign layer_1_weights[11][19] = 6'sd6;
    assign layer_1_weights[11][20] = 6'sd5;
    assign layer_1_weights[11][21] = -6'sd3;
    assign layer_1_weights[11][22] = -6'sd4;
    assign layer_1_weights[11][23] = 6'sd3;
    assign layer_1_weights[11][24] = -6'sd1;
    assign layer_1_weights[11][25] = -6'sd3;
    assign layer_1_weights[11][26] = -6'sd8;
    assign layer_1_weights[11][27] = -6'sd2;
    assign layer_1_weights[11][28] = -6'sd6;
    assign layer_1_weights[11][29] = -6'sd6;
    assign layer_1_weights[11][30] = 6'sd2;
    assign layer_1_weights[11][31] = 6'sd6;
    assign layer_1_weights[11][32] = 6'sd2;
    assign layer_1_weights[11][33] = -6'sd3;
    assign layer_1_weights[11][34] = -6'sd2;
    assign layer_1_weights[11][35] = 6'sd1;
    assign layer_1_weights[11][36] = -6'sd1;
    assign layer_1_weights[11][37] = -6'sd4;
    assign layer_1_weights[11][38] = -6'sd9;
    assign layer_1_weights[11][39] = -6'sd7;
    assign layer_1_weights[11][40] = -6'sd2;
    assign layer_1_weights[11][41] = 6'sd1;
    assign layer_1_weights[11][42] = 6'sd1;
    assign layer_1_weights[11][43] = 6'sd1;
    assign layer_1_weights[11][44] = 6'sd2;
    assign layer_1_weights[11][45] = 6'sd1;
    assign layer_1_weights[11][46] = -6'sd2;
    assign layer_1_weights[11][47] = -6'sd1;
    assign layer_1_weights[11][48] = 6'sd0;
    assign layer_1_weights[11][49] = -6'sd5;
    assign layer_1_weights[11][50] = -6'sd4;
    assign layer_1_weights[11][51] = -6'sd1;
    assign layer_1_weights[11][52] = 6'sd1;
    assign layer_1_weights[11][53] = 6'sd0;
    assign layer_1_weights[11][54] = -6'sd2;
    assign layer_1_weights[11][55] = -6'sd1;
    assign layer_1_weights[11][56] = 6'sd3;
    assign layer_1_weights[11][57] = 6'sd3;
    assign layer_1_weights[11][58] = -6'sd2;
    assign layer_1_weights[11][59] = -6'sd1;
    assign layer_1_weights[11][60] = -6'sd5;
    assign layer_1_weights[11][61] = 6'sd3;
    assign layer_1_weights[11][62] = -6'sd1;
    assign layer_1_weights[11][63] = 6'sd1;
    assign layer_1_weights[11][64] = -6'sd3;
    assign layer_1_weights[11][65] = 6'sd0;
    assign layer_1_weights[11][66] = 6'sd2;
    assign layer_1_weights[11][67] = 6'sd2;
    assign layer_1_weights[11][68] = 6'sd3;
    assign layer_1_weights[11][69] = 6'sd1;
    assign layer_1_weights[11][70] = -6'sd2;
    assign layer_1_weights[11][71] = 6'sd0;
    assign layer_1_weights[11][72] = -6'sd3;
    assign layer_1_weights[11][73] = -6'sd2;
    assign layer_1_weights[11][74] = 6'sd0;
    assign layer_1_weights[11][75] = -6'sd1;
    assign layer_1_weights[11][76] = -6'sd1;
    assign layer_1_weights[11][77] = 6'sd4;
    assign layer_1_weights[11][78] = 6'sd7;
    assign layer_1_weights[11][79] = -6'sd1;
    assign layer_1_weights[11][80] = -6'sd5;
    assign layer_1_weights[11][81] = -6'sd1;
    assign layer_1_weights[11][82] = -6'sd2;
    assign layer_1_weights[11][83] = 6'sd7;
    assign layer_1_weights[11][84] = -6'sd3;
    assign layer_1_weights[11][85] = 6'sd1;
    assign layer_1_weights[11][86] = -6'sd2;
    assign layer_1_weights[11][87] = 6'sd2;
    assign layer_1_weights[11][88] = 6'sd2;
    assign layer_1_weights[11][89] = 6'sd2;
    assign layer_1_weights[11][90] = 6'sd0;
    assign layer_1_weights[11][91] = -6'sd6;
    assign layer_1_weights[11][92] = -6'sd8;
    assign layer_1_weights[11][93] = -6'sd2;
    assign layer_1_weights[11][94] = 6'sd2;
    assign layer_1_weights[11][95] = 6'sd3;
    assign layer_1_weights[11][96] = -6'sd3;
    assign layer_1_weights[11][97] = -6'sd3;
    assign layer_1_weights[11][98] = 6'sd0;
    assign layer_1_weights[11][99] = 6'sd2;
    assign layer_1_weights[11][100] = 6'sd3;
    assign layer_1_weights[11][101] = 6'sd2;
    assign layer_1_weights[11][102] = 6'sd1;
    assign layer_1_weights[11][103] = 6'sd2;
    assign layer_1_weights[11][104] = 6'sd1;
    assign layer_1_weights[11][105] = 6'sd4;
    assign layer_1_weights[11][106] = 6'sd7;
    assign layer_1_weights[11][107] = 6'sd10;
    assign layer_1_weights[11][108] = 6'sd2;
    assign layer_1_weights[11][109] = 6'sd5;
    assign layer_1_weights[11][110] = 6'sd3;
    assign layer_1_weights[11][111] = 6'sd2;
    assign layer_1_weights[11][112] = -6'sd1;
    assign layer_1_weights[11][113] = 6'sd2;
    assign layer_1_weights[11][114] = 6'sd4;
    assign layer_1_weights[11][115] = 6'sd3;
    assign layer_1_weights[11][116] = 6'sd5;
    assign layer_1_weights[11][117] = 6'sd0;
    assign layer_1_weights[11][118] = 6'sd2;
    assign layer_1_weights[11][119] = -6'sd3;
    assign layer_1_weights[11][120] = -6'sd1;
    assign layer_1_weights[11][121] = -6'sd2;
    assign layer_1_weights[11][122] = 6'sd2;
    assign layer_1_weights[11][123] = 6'sd0;
    assign layer_1_weights[11][124] = -6'sd1;
    assign layer_1_weights[11][125] = 6'sd0;
    assign layer_1_weights[11][126] = 6'sd0;
    assign layer_1_weights[11][127] = 6'sd1;
    assign layer_1_weights[11][128] = 6'sd2;
    assign layer_1_weights[11][129] = 6'sd3;
    assign layer_1_weights[11][130] = 6'sd0;
    assign layer_1_weights[11][131] = 6'sd8;
    assign layer_1_weights[11][132] = 6'sd0;
    assign layer_1_weights[11][133] = 6'sd1;
    assign layer_1_weights[11][134] = -6'sd1;
    assign layer_1_weights[11][135] = 6'sd2;
    assign layer_1_weights[11][136] = -6'sd1;
    assign layer_1_weights[11][137] = 6'sd3;
    assign layer_1_weights[11][138] = 6'sd3;
    assign layer_1_weights[11][139] = 6'sd7;
    assign layer_1_weights[11][140] = 6'sd0;
    assign layer_1_weights[11][141] = 6'sd0;
    assign layer_1_weights[11][142] = -6'sd1;
    assign layer_1_weights[11][143] = -6'sd1;
    assign layer_1_biases[11] = -6'sd1;
    assign layer_1_weights[12][0] = 6'sd2;
    assign layer_1_weights[12][1] = -6'sd1;
    assign layer_1_weights[12][2] = -6'sd2;
    assign layer_1_weights[12][3] = -6'sd2;
    assign layer_1_weights[12][4] = -6'sd5;
    assign layer_1_weights[12][5] = -6'sd10;
    assign layer_1_weights[12][6] = 6'sd0;
    assign layer_1_weights[12][7] = 6'sd8;
    assign layer_1_weights[12][8] = 6'sd1;
    assign layer_1_weights[12][9] = 6'sd7;
    assign layer_1_weights[12][10] = -6'sd1;
    assign layer_1_weights[12][11] = -6'sd1;
    assign layer_1_weights[12][12] = 6'sd0;
    assign layer_1_weights[12][13] = 6'sd0;
    assign layer_1_weights[12][14] = 6'sd0;
    assign layer_1_weights[12][15] = 6'sd3;
    assign layer_1_weights[12][16] = 6'sd3;
    assign layer_1_weights[12][17] = 6'sd2;
    assign layer_1_weights[12][18] = -6'sd2;
    assign layer_1_weights[12][19] = 6'sd1;
    assign layer_1_weights[12][20] = 6'sd4;
    assign layer_1_weights[12][21] = 6'sd4;
    assign layer_1_weights[12][22] = 6'sd3;
    assign layer_1_weights[12][23] = 6'sd5;
    assign layer_1_weights[12][24] = 6'sd1;
    assign layer_1_weights[12][25] = -6'sd4;
    assign layer_1_weights[12][26] = -6'sd8;
    assign layer_1_weights[12][27] = -6'sd2;
    assign layer_1_weights[12][28] = -6'sd5;
    assign layer_1_weights[12][29] = -6'sd4;
    assign layer_1_weights[12][30] = 6'sd0;
    assign layer_1_weights[12][31] = 6'sd3;
    assign layer_1_weights[12][32] = 6'sd5;
    assign layer_1_weights[12][33] = 6'sd2;
    assign layer_1_weights[12][34] = 6'sd5;
    assign layer_1_weights[12][35] = 6'sd8;
    assign layer_1_weights[12][36] = 6'sd4;
    assign layer_1_weights[12][37] = -6'sd9;
    assign layer_1_weights[12][38] = -6'sd5;
    assign layer_1_weights[12][39] = -6'sd5;
    assign layer_1_weights[12][40] = -6'sd3;
    assign layer_1_weights[12][41] = -6'sd2;
    assign layer_1_weights[12][42] = 6'sd4;
    assign layer_1_weights[12][43] = 6'sd2;
    assign layer_1_weights[12][44] = 6'sd2;
    assign layer_1_weights[12][45] = 6'sd1;
    assign layer_1_weights[12][46] = -6'sd1;
    assign layer_1_weights[12][47] = 6'sd10;
    assign layer_1_weights[12][48] = -6'sd4;
    assign layer_1_weights[12][49] = -6'sd8;
    assign layer_1_weights[12][50] = 6'sd2;
    assign layer_1_weights[12][51] = -6'sd2;
    assign layer_1_weights[12][52] = -6'sd2;
    assign layer_1_weights[12][53] = 6'sd4;
    assign layer_1_weights[12][54] = 6'sd0;
    assign layer_1_weights[12][55] = -6'sd2;
    assign layer_1_weights[12][56] = -6'sd1;
    assign layer_1_weights[12][57] = -6'sd2;
    assign layer_1_weights[12][58] = -6'sd2;
    assign layer_1_weights[12][59] = -6'sd1;
    assign layer_1_weights[12][60] = -6'sd1;
    assign layer_1_weights[12][61] = -6'sd5;
    assign layer_1_weights[12][62] = -6'sd8;
    assign layer_1_weights[12][63] = -6'sd6;
    assign layer_1_weights[12][64] = -6'sd2;
    assign layer_1_weights[12][65] = 6'sd6;
    assign layer_1_weights[12][66] = 6'sd4;
    assign layer_1_weights[12][67] = -6'sd3;
    assign layer_1_weights[12][68] = 6'sd1;
    assign layer_1_weights[12][69] = -6'sd3;
    assign layer_1_weights[12][70] = -6'sd4;
    assign layer_1_weights[12][71] = 6'sd6;
    assign layer_1_weights[12][72] = -6'sd2;
    assign layer_1_weights[12][73] = 6'sd0;
    assign layer_1_weights[12][74] = -6'sd2;
    assign layer_1_weights[12][75] = -6'sd4;
    assign layer_1_weights[12][76] = -6'sd2;
    assign layer_1_weights[12][77] = 6'sd3;
    assign layer_1_weights[12][78] = -6'sd2;
    assign layer_1_weights[12][79] = 6'sd0;
    assign layer_1_weights[12][80] = -6'sd1;
    assign layer_1_weights[12][81] = -6'sd3;
    assign layer_1_weights[12][82] = -6'sd8;
    assign layer_1_weights[12][83] = -6'sd6;
    assign layer_1_weights[12][84] = 6'sd5;
    assign layer_1_weights[12][85] = 6'sd5;
    assign layer_1_weights[12][86] = 6'sd3;
    assign layer_1_weights[12][87] = -6'sd1;
    assign layer_1_weights[12][88] = -6'sd4;
    assign layer_1_weights[12][89] = -6'sd3;
    assign layer_1_weights[12][90] = 6'sd1;
    assign layer_1_weights[12][91] = 6'sd6;
    assign layer_1_weights[12][92] = 6'sd0;
    assign layer_1_weights[12][93] = -6'sd6;
    assign layer_1_weights[12][94] = -6'sd9;
    assign layer_1_weights[12][95] = -6'sd3;
    assign layer_1_weights[12][96] = 6'sd4;
    assign layer_1_weights[12][97] = 6'sd3;
    assign layer_1_weights[12][98] = 6'sd3;
    assign layer_1_weights[12][99] = 6'sd1;
    assign layer_1_weights[12][100] = 6'sd1;
    assign layer_1_weights[12][101] = -6'sd2;
    assign layer_1_weights[12][102] = 6'sd2;
    assign layer_1_weights[12][103] = 6'sd8;
    assign layer_1_weights[12][104] = -6'sd2;
    assign layer_1_weights[12][105] = -6'sd10;
    assign layer_1_weights[12][106] = -6'sd12;
    assign layer_1_weights[12][107] = 6'sd4;
    assign layer_1_weights[12][108] = -6'sd2;
    assign layer_1_weights[12][109] = -6'sd2;
    assign layer_1_weights[12][110] = 6'sd2;
    assign layer_1_weights[12][111] = 6'sd1;
    assign layer_1_weights[12][112] = 6'sd5;
    assign layer_1_weights[12][113] = 6'sd5;
    assign layer_1_weights[12][114] = 6'sd4;
    assign layer_1_weights[12][115] = 6'sd2;
    assign layer_1_weights[12][116] = -6'sd7;
    assign layer_1_weights[12][117] = -6'sd8;
    assign layer_1_weights[12][118] = -6'sd11;
    assign layer_1_weights[12][119] = 6'sd1;
    assign layer_1_weights[12][120] = 6'sd0;
    assign layer_1_weights[12][121] = -6'sd1;
    assign layer_1_weights[12][122] = 6'sd1;
    assign layer_1_weights[12][123] = 6'sd2;
    assign layer_1_weights[12][124] = 6'sd1;
    assign layer_1_weights[12][125] = 6'sd4;
    assign layer_1_weights[12][126] = 6'sd2;
    assign layer_1_weights[12][127] = -6'sd6;
    assign layer_1_weights[12][128] = -6'sd10;
    assign layer_1_weights[12][129] = -6'sd9;
    assign layer_1_weights[12][130] = -6'sd7;
    assign layer_1_weights[12][131] = 6'sd1;
    assign layer_1_weights[12][132] = 6'sd2;
    assign layer_1_weights[12][133] = 6'sd5;
    assign layer_1_weights[12][134] = -6'sd2;
    assign layer_1_weights[12][135] = -6'sd3;
    assign layer_1_weights[12][136] = -6'sd9;
    assign layer_1_weights[12][137] = -6'sd6;
    assign layer_1_weights[12][138] = -6'sd2;
    assign layer_1_weights[12][139] = 6'sd7;
    assign layer_1_weights[12][140] = -6'sd4;
    assign layer_1_weights[12][141] = 6'sd6;
    assign layer_1_weights[12][142] = -6'sd1;
    assign layer_1_weights[12][143] = 6'sd1;
    assign layer_1_biases[12] = -6'sd6;
    assign layer_1_weights[13][0] = 6'sd0;
    assign layer_1_weights[13][1] = 6'sd1;
    assign layer_1_weights[13][2] = -6'sd2;
    assign layer_1_weights[13][3] = -6'sd4;
    assign layer_1_weights[13][4] = 6'sd2;
    assign layer_1_weights[13][5] = -6'sd5;
    assign layer_1_weights[13][6] = 6'sd0;
    assign layer_1_weights[13][7] = 6'sd0;
    assign layer_1_weights[13][8] = -6'sd3;
    assign layer_1_weights[13][9] = -6'sd3;
    assign layer_1_weights[13][10] = -6'sd2;
    assign layer_1_weights[13][11] = 6'sd1;
    assign layer_1_weights[13][12] = -6'sd1;
    assign layer_1_weights[13][13] = 6'sd1;
    assign layer_1_weights[13][14] = 6'sd2;
    assign layer_1_weights[13][15] = 6'sd5;
    assign layer_1_weights[13][16] = 6'sd3;
    assign layer_1_weights[13][17] = 6'sd1;
    assign layer_1_weights[13][18] = 6'sd1;
    assign layer_1_weights[13][19] = 6'sd2;
    assign layer_1_weights[13][20] = -6'sd3;
    assign layer_1_weights[13][21] = 6'sd0;
    assign layer_1_weights[13][22] = -6'sd8;
    assign layer_1_weights[13][23] = 6'sd1;
    assign layer_1_weights[13][24] = 6'sd1;
    assign layer_1_weights[13][25] = -6'sd1;
    assign layer_1_weights[13][26] = 6'sd5;
    assign layer_1_weights[13][27] = 6'sd2;
    assign layer_1_weights[13][28] = 6'sd4;
    assign layer_1_weights[13][29] = 6'sd5;
    assign layer_1_weights[13][30] = 6'sd3;
    assign layer_1_weights[13][31] = -6'sd2;
    assign layer_1_weights[13][32] = 6'sd3;
    assign layer_1_weights[13][33] = -6'sd2;
    assign layer_1_weights[13][34] = -6'sd6;
    assign layer_1_weights[13][35] = -6'sd2;
    assign layer_1_weights[13][36] = 6'sd5;
    assign layer_1_weights[13][37] = 6'sd13;
    assign layer_1_weights[13][38] = 6'sd8;
    assign layer_1_weights[13][39] = 6'sd5;
    assign layer_1_weights[13][40] = 6'sd5;
    assign layer_1_weights[13][41] = 6'sd4;
    assign layer_1_weights[13][42] = -6'sd2;
    assign layer_1_weights[13][43] = -6'sd1;
    assign layer_1_weights[13][44] = 6'sd4;
    assign layer_1_weights[13][45] = 6'sd1;
    assign layer_1_weights[13][46] = -6'sd2;
    assign layer_1_weights[13][47] = -6'sd6;
    assign layer_1_weights[13][48] = 6'sd0;
    assign layer_1_weights[13][49] = -6'sd6;
    assign layer_1_weights[13][50] = -6'sd8;
    assign layer_1_weights[13][51] = -6'sd8;
    assign layer_1_weights[13][52] = -6'sd9;
    assign layer_1_weights[13][53] = -6'sd2;
    assign layer_1_weights[13][54] = -6'sd1;
    assign layer_1_weights[13][55] = 6'sd1;
    assign layer_1_weights[13][56] = 6'sd3;
    assign layer_1_weights[13][57] = -6'sd1;
    assign layer_1_weights[13][58] = 6'sd1;
    assign layer_1_weights[13][59] = 6'sd3;
    assign layer_1_weights[13][60] = -6'sd2;
    assign layer_1_weights[13][61] = -6'sd18;
    assign layer_1_weights[13][62] = -6'sd13;
    assign layer_1_weights[13][63] = -6'sd9;
    assign layer_1_weights[13][64] = -6'sd4;
    assign layer_1_weights[13][65] = 6'sd3;
    assign layer_1_weights[13][66] = -6'sd1;
    assign layer_1_weights[13][67] = 6'sd1;
    assign layer_1_weights[13][68] = -6'sd2;
    assign layer_1_weights[13][69] = -6'sd2;
    assign layer_1_weights[13][70] = -6'sd1;
    assign layer_1_weights[13][71] = -6'sd4;
    assign layer_1_weights[13][72] = 6'sd2;
    assign layer_1_weights[13][73] = 6'sd6;
    assign layer_1_weights[13][74] = 6'sd4;
    assign layer_1_weights[13][75] = 6'sd4;
    assign layer_1_weights[13][76] = 6'sd7;
    assign layer_1_weights[13][77] = 6'sd3;
    assign layer_1_weights[13][78] = -6'sd1;
    assign layer_1_weights[13][79] = -6'sd1;
    assign layer_1_weights[13][80] = 6'sd0;
    assign layer_1_weights[13][81] = 6'sd4;
    assign layer_1_weights[13][82] = 6'sd4;
    assign layer_1_weights[13][83] = 6'sd0;
    assign layer_1_weights[13][84] = 6'sd7;
    assign layer_1_weights[13][85] = 6'sd6;
    assign layer_1_weights[13][86] = 6'sd5;
    assign layer_1_weights[13][87] = 6'sd2;
    assign layer_1_weights[13][88] = 6'sd3;
    assign layer_1_weights[13][89] = -6'sd4;
    assign layer_1_weights[13][90] = 6'sd2;
    assign layer_1_weights[13][91] = -6'sd1;
    assign layer_1_weights[13][92] = -6'sd1;
    assign layer_1_weights[13][93] = 6'sd3;
    assign layer_1_weights[13][94] = 6'sd2;
    assign layer_1_weights[13][95] = 6'sd0;
    assign layer_1_weights[13][96] = -6'sd1;
    assign layer_1_weights[13][97] = 6'sd3;
    assign layer_1_weights[13][98] = 6'sd2;
    assign layer_1_weights[13][99] = 6'sd2;
    assign layer_1_weights[13][100] = 6'sd0;
    assign layer_1_weights[13][101] = -6'sd4;
    assign layer_1_weights[13][102] = 6'sd0;
    assign layer_1_weights[13][103] = -6'sd2;
    assign layer_1_weights[13][104] = -6'sd2;
    assign layer_1_weights[13][105] = -6'sd2;
    assign layer_1_weights[13][106] = 6'sd1;
    assign layer_1_weights[13][107] = -6'sd2;
    assign layer_1_weights[13][108] = 6'sd6;
    assign layer_1_weights[13][109] = 6'sd2;
    assign layer_1_weights[13][110] = 6'sd0;
    assign layer_1_weights[13][111] = 6'sd0;
    assign layer_1_weights[13][112] = 6'sd0;
    assign layer_1_weights[13][113] = 6'sd0;
    assign layer_1_weights[13][114] = -6'sd1;
    assign layer_1_weights[13][115] = -6'sd4;
    assign layer_1_weights[13][116] = 6'sd2;
    assign layer_1_weights[13][117] = -6'sd3;
    assign layer_1_weights[13][118] = 6'sd0;
    assign layer_1_weights[13][119] = 6'sd2;
    assign layer_1_weights[13][120] = -6'sd1;
    assign layer_1_weights[13][121] = 6'sd3;
    assign layer_1_weights[13][122] = 6'sd3;
    assign layer_1_weights[13][123] = 6'sd4;
    assign layer_1_weights[13][124] = 6'sd2;
    assign layer_1_weights[13][125] = 6'sd2;
    assign layer_1_weights[13][126] = 6'sd1;
    assign layer_1_weights[13][127] = 6'sd1;
    assign layer_1_weights[13][128] = -6'sd3;
    assign layer_1_weights[13][129] = -6'sd4;
    assign layer_1_weights[13][130] = -6'sd2;
    assign layer_1_weights[13][131] = 6'sd1;
    assign layer_1_weights[13][132] = 6'sd0;
    assign layer_1_weights[13][133] = -6'sd6;
    assign layer_1_weights[13][134] = 6'sd0;
    assign layer_1_weights[13][135] = 6'sd5;
    assign layer_1_weights[13][136] = 6'sd6;
    assign layer_1_weights[13][137] = 6'sd7;
    assign layer_1_weights[13][138] = 6'sd7;
    assign layer_1_weights[13][139] = 6'sd13;
    assign layer_1_weights[13][140] = 6'sd9;
    assign layer_1_weights[13][141] = 6'sd7;
    assign layer_1_weights[13][142] = 6'sd2;
    assign layer_1_weights[13][143] = 6'sd0;
    assign layer_1_biases[13] = -6'sd3;
    assign layer_1_weights[14][0] = 6'sd0;
    assign layer_1_weights[14][1] = -6'sd1;
    assign layer_1_weights[14][2] = -6'sd3;
    assign layer_1_weights[14][3] = -6'sd9;
    assign layer_1_weights[14][4] = -6'sd4;
    assign layer_1_weights[14][5] = -6'sd5;
    assign layer_1_weights[14][6] = -6'sd11;
    assign layer_1_weights[14][7] = -6'sd1;
    assign layer_1_weights[14][8] = -6'sd4;
    assign layer_1_weights[14][9] = -6'sd6;
    assign layer_1_weights[14][10] = 6'sd1;
    assign layer_1_weights[14][11] = 6'sd0;
    assign layer_1_weights[14][12] = 6'sd1;
    assign layer_1_weights[14][13] = 6'sd1;
    assign layer_1_weights[14][14] = -6'sd6;
    assign layer_1_weights[14][15] = -6'sd1;
    assign layer_1_weights[14][16] = 6'sd0;
    assign layer_1_weights[14][17] = -6'sd2;
    assign layer_1_weights[14][18] = 6'sd2;
    assign layer_1_weights[14][19] = 6'sd3;
    assign layer_1_weights[14][20] = 6'sd2;
    assign layer_1_weights[14][21] = 6'sd5;
    assign layer_1_weights[14][22] = -6'sd2;
    assign layer_1_weights[14][23] = 6'sd1;
    assign layer_1_weights[14][24] = -6'sd1;
    assign layer_1_weights[14][25] = 6'sd1;
    assign layer_1_weights[14][26] = 6'sd10;
    assign layer_1_weights[14][27] = 6'sd3;
    assign layer_1_weights[14][28] = 6'sd1;
    assign layer_1_weights[14][29] = -6'sd5;
    assign layer_1_weights[14][30] = -6'sd1;
    assign layer_1_weights[14][31] = 6'sd7;
    assign layer_1_weights[14][32] = 6'sd4;
    assign layer_1_weights[14][33] = 6'sd0;
    assign layer_1_weights[14][34] = -6'sd3;
    assign layer_1_weights[14][35] = 6'sd4;
    assign layer_1_weights[14][36] = 6'sd2;
    assign layer_1_weights[14][37] = 6'sd0;
    assign layer_1_weights[14][38] = 6'sd6;
    assign layer_1_weights[14][39] = 6'sd3;
    assign layer_1_weights[14][40] = 6'sd0;
    assign layer_1_weights[14][41] = -6'sd6;
    assign layer_1_weights[14][42] = 6'sd1;
    assign layer_1_weights[14][43] = 6'sd9;
    assign layer_1_weights[14][44] = -6'sd2;
    assign layer_1_weights[14][45] = -6'sd5;
    assign layer_1_weights[14][46] = 6'sd2;
    assign layer_1_weights[14][47] = 6'sd8;
    assign layer_1_weights[14][48] = 6'sd7;
    assign layer_1_weights[14][49] = 6'sd0;
    assign layer_1_weights[14][50] = -6'sd1;
    assign layer_1_weights[14][51] = 6'sd3;
    assign layer_1_weights[14][52] = 6'sd1;
    assign layer_1_weights[14][53] = -6'sd3;
    assign layer_1_weights[14][54] = 6'sd2;
    assign layer_1_weights[14][55] = 6'sd3;
    assign layer_1_weights[14][56] = -6'sd3;
    assign layer_1_weights[14][57] = -6'sd5;
    assign layer_1_weights[14][58] = -6'sd14;
    assign layer_1_weights[14][59] = -6'sd5;
    assign layer_1_weights[14][60] = 6'sd3;
    assign layer_1_weights[14][61] = -6'sd2;
    assign layer_1_weights[14][62] = -6'sd2;
    assign layer_1_weights[14][63] = 6'sd0;
    assign layer_1_weights[14][64] = 6'sd0;
    assign layer_1_weights[14][65] = -6'sd3;
    assign layer_1_weights[14][66] = 6'sd0;
    assign layer_1_weights[14][67] = -6'sd3;
    assign layer_1_weights[14][68] = -6'sd5;
    assign layer_1_weights[14][69] = -6'sd3;
    assign layer_1_weights[14][70] = -6'sd2;
    assign layer_1_weights[14][71] = 6'sd1;
    assign layer_1_weights[14][72] = 6'sd3;
    assign layer_1_weights[14][73] = -6'sd1;
    assign layer_1_weights[14][74] = 6'sd0;
    assign layer_1_weights[14][75] = 6'sd1;
    assign layer_1_weights[14][76] = 6'sd1;
    assign layer_1_weights[14][77] = -6'sd1;
    assign layer_1_weights[14][78] = -6'sd1;
    assign layer_1_weights[14][79] = 6'sd0;
    assign layer_1_weights[14][80] = -6'sd1;
    assign layer_1_weights[14][81] = 6'sd7;
    assign layer_1_weights[14][82] = 6'sd6;
    assign layer_1_weights[14][83] = 6'sd5;
    assign layer_1_weights[14][84] = -6'sd4;
    assign layer_1_weights[14][85] = 6'sd3;
    assign layer_1_weights[14][86] = 6'sd3;
    assign layer_1_weights[14][87] = 6'sd2;
    assign layer_1_weights[14][88] = -6'sd3;
    assign layer_1_weights[14][89] = -6'sd2;
    assign layer_1_weights[14][90] = 6'sd2;
    assign layer_1_weights[14][91] = 6'sd1;
    assign layer_1_weights[14][92] = 6'sd1;
    assign layer_1_weights[14][93] = 6'sd4;
    assign layer_1_weights[14][94] = 6'sd5;
    assign layer_1_weights[14][95] = 6'sd3;
    assign layer_1_weights[14][96] = -6'sd5;
    assign layer_1_weights[14][97] = 6'sd6;
    assign layer_1_weights[14][98] = 6'sd1;
    assign layer_1_weights[14][99] = 6'sd1;
    assign layer_1_weights[14][100] = -6'sd8;
    assign layer_1_weights[14][101] = -6'sd2;
    assign layer_1_weights[14][102] = 6'sd3;
    assign layer_1_weights[14][103] = 6'sd3;
    assign layer_1_weights[14][104] = -6'sd1;
    assign layer_1_weights[14][105] = 6'sd5;
    assign layer_1_weights[14][106] = 6'sd2;
    assign layer_1_weights[14][107] = -6'sd4;
    assign layer_1_weights[14][108] = 6'sd5;
    assign layer_1_weights[14][109] = 6'sd0;
    assign layer_1_weights[14][110] = 6'sd1;
    assign layer_1_weights[14][111] = -6'sd1;
    assign layer_1_weights[14][112] = -6'sd1;
    assign layer_1_weights[14][113] = 6'sd3;
    assign layer_1_weights[14][114] = 6'sd0;
    assign layer_1_weights[14][115] = 6'sd0;
    assign layer_1_weights[14][116] = 6'sd3;
    assign layer_1_weights[14][117] = 6'sd4;
    assign layer_1_weights[14][118] = 6'sd3;
    assign layer_1_weights[14][119] = 6'sd2;
    assign layer_1_weights[14][120] = 6'sd0;
    assign layer_1_weights[14][121] = 6'sd11;
    assign layer_1_weights[14][122] = 6'sd3;
    assign layer_1_weights[14][123] = 6'sd2;
    assign layer_1_weights[14][124] = -6'sd5;
    assign layer_1_weights[14][125] = -6'sd4;
    assign layer_1_weights[14][126] = -6'sd2;
    assign layer_1_weights[14][127] = 6'sd1;
    assign layer_1_weights[14][128] = 6'sd0;
    assign layer_1_weights[14][129] = -6'sd3;
    assign layer_1_weights[14][130] = 6'sd0;
    assign layer_1_weights[14][131] = 6'sd6;
    assign layer_1_weights[14][132] = -6'sd2;
    assign layer_1_weights[14][133] = -6'sd2;
    assign layer_1_weights[14][134] = -6'sd6;
    assign layer_1_weights[14][135] = 6'sd6;
    assign layer_1_weights[14][136] = 6'sd1;
    assign layer_1_weights[14][137] = -6'sd2;
    assign layer_1_weights[14][138] = -6'sd2;
    assign layer_1_weights[14][139] = 6'sd0;
    assign layer_1_weights[14][140] = -6'sd4;
    assign layer_1_weights[14][141] = 6'sd4;
    assign layer_1_weights[14][142] = 6'sd1;
    assign layer_1_weights[14][143] = 6'sd0;
    assign layer_1_biases[14] = 6'sd3;
    assign layer_1_weights[15][0] = 6'sd1;
    assign layer_1_weights[15][1] = -6'sd2;
    assign layer_1_weights[15][2] = -6'sd2;
    assign layer_1_weights[15][3] = 6'sd4;
    assign layer_1_weights[15][4] = 6'sd7;
    assign layer_1_weights[15][5] = 6'sd2;
    assign layer_1_weights[15][6] = 6'sd0;
    assign layer_1_weights[15][7] = 6'sd0;
    assign layer_1_weights[15][8] = 6'sd3;
    assign layer_1_weights[15][9] = -6'sd2;
    assign layer_1_weights[15][10] = 6'sd1;
    assign layer_1_weights[15][11] = 6'sd0;
    assign layer_1_weights[15][12] = 6'sd1;
    assign layer_1_weights[15][13] = 6'sd0;
    assign layer_1_weights[15][14] = 6'sd3;
    assign layer_1_weights[15][15] = 6'sd5;
    assign layer_1_weights[15][16] = 6'sd3;
    assign layer_1_weights[15][17] = 6'sd3;
    assign layer_1_weights[15][18] = 6'sd0;
    assign layer_1_weights[15][19] = -6'sd1;
    assign layer_1_weights[15][20] = -6'sd2;
    assign layer_1_weights[15][21] = -6'sd2;
    assign layer_1_weights[15][22] = -6'sd1;
    assign layer_1_weights[15][23] = 6'sd3;
    assign layer_1_weights[15][24] = 6'sd0;
    assign layer_1_weights[15][25] = -6'sd7;
    assign layer_1_weights[15][26] = 6'sd6;
    assign layer_1_weights[15][27] = 6'sd4;
    assign layer_1_weights[15][28] = 6'sd4;
    assign layer_1_weights[15][29] = 6'sd4;
    assign layer_1_weights[15][30] = 6'sd10;
    assign layer_1_weights[15][31] = 6'sd10;
    assign layer_1_weights[15][32] = 6'sd3;
    assign layer_1_weights[15][33] = 6'sd4;
    assign layer_1_weights[15][34] = -6'sd2;
    assign layer_1_weights[15][35] = 6'sd0;
    assign layer_1_weights[15][36] = -6'sd2;
    assign layer_1_weights[15][37] = 6'sd4;
    assign layer_1_weights[15][38] = 6'sd4;
    assign layer_1_weights[15][39] = 6'sd1;
    assign layer_1_weights[15][40] = 6'sd4;
    assign layer_1_weights[15][41] = 6'sd4;
    assign layer_1_weights[15][42] = 6'sd7;
    assign layer_1_weights[15][43] = 6'sd9;
    assign layer_1_weights[15][44] = 6'sd6;
    assign layer_1_weights[15][45] = 6'sd3;
    assign layer_1_weights[15][46] = 6'sd4;
    assign layer_1_weights[15][47] = 6'sd2;
    assign layer_1_weights[15][48] = -6'sd4;
    assign layer_1_weights[15][49] = -6'sd4;
    assign layer_1_weights[15][50] = -6'sd3;
    assign layer_1_weights[15][51] = -6'sd6;
    assign layer_1_weights[15][52] = -6'sd3;
    assign layer_1_weights[15][53] = -6'sd8;
    assign layer_1_weights[15][54] = -6'sd8;
    assign layer_1_weights[15][55] = -6'sd1;
    assign layer_1_weights[15][56] = -6'sd1;
    assign layer_1_weights[15][57] = 6'sd0;
    assign layer_1_weights[15][58] = -6'sd3;
    assign layer_1_weights[15][59] = 6'sd4;
    assign layer_1_weights[15][60] = -6'sd5;
    assign layer_1_weights[15][61] = -6'sd8;
    assign layer_1_weights[15][62] = -6'sd3;
    assign layer_1_weights[15][63] = -6'sd3;
    assign layer_1_weights[15][64] = -6'sd4;
    assign layer_1_weights[15][65] = -6'sd3;
    assign layer_1_weights[15][66] = -6'sd3;
    assign layer_1_weights[15][67] = -6'sd3;
    assign layer_1_weights[15][68] = 6'sd2;
    assign layer_1_weights[15][69] = -6'sd1;
    assign layer_1_weights[15][70] = -6'sd6;
    assign layer_1_weights[15][71] = -6'sd4;
    assign layer_1_weights[15][72] = -6'sd4;
    assign layer_1_weights[15][73] = 6'sd0;
    assign layer_1_weights[15][74] = 6'sd4;
    assign layer_1_weights[15][75] = 6'sd1;
    assign layer_1_weights[15][76] = -6'sd1;
    assign layer_1_weights[15][77] = 6'sd3;
    assign layer_1_weights[15][78] = -6'sd1;
    assign layer_1_weights[15][79] = -6'sd1;
    assign layer_1_weights[15][80] = 6'sd0;
    assign layer_1_weights[15][81] = 6'sd1;
    assign layer_1_weights[15][82] = -6'sd1;
    assign layer_1_weights[15][83] = 6'sd3;
    assign layer_1_weights[15][84] = -6'sd5;
    assign layer_1_weights[15][85] = 6'sd4;
    assign layer_1_weights[15][86] = 6'sd1;
    assign layer_1_weights[15][87] = 6'sd1;
    assign layer_1_weights[15][88] = 6'sd0;
    assign layer_1_weights[15][89] = -6'sd2;
    assign layer_1_weights[15][90] = -6'sd2;
    assign layer_1_weights[15][91] = 6'sd1;
    assign layer_1_weights[15][92] = -6'sd4;
    assign layer_1_weights[15][93] = -6'sd2;
    assign layer_1_weights[15][94] = -6'sd3;
    assign layer_1_weights[15][95] = -6'sd1;
    assign layer_1_weights[15][96] = 6'sd7;
    assign layer_1_weights[15][97] = 6'sd1;
    assign layer_1_weights[15][98] = -6'sd1;
    assign layer_1_weights[15][99] = 6'sd4;
    assign layer_1_weights[15][100] = -6'sd1;
    assign layer_1_weights[15][101] = -6'sd2;
    assign layer_1_weights[15][102] = 6'sd3;
    assign layer_1_weights[15][103] = 6'sd2;
    assign layer_1_weights[15][104] = -6'sd1;
    assign layer_1_weights[15][105] = -6'sd3;
    assign layer_1_weights[15][106] = 6'sd2;
    assign layer_1_weights[15][107] = 6'sd2;
    assign layer_1_weights[15][108] = 6'sd5;
    assign layer_1_weights[15][109] = 6'sd0;
    assign layer_1_weights[15][110] = 6'sd3;
    assign layer_1_weights[15][111] = 6'sd3;
    assign layer_1_weights[15][112] = 6'sd4;
    assign layer_1_weights[15][113] = 6'sd4;
    assign layer_1_weights[15][114] = 6'sd1;
    assign layer_1_weights[15][115] = -6'sd3;
    assign layer_1_weights[15][116] = 6'sd1;
    assign layer_1_weights[15][117] = 6'sd0;
    assign layer_1_weights[15][118] = 6'sd6;
    assign layer_1_weights[15][119] = 6'sd3;
    assign layer_1_weights[15][120] = 6'sd1;
    assign layer_1_weights[15][121] = 6'sd6;
    assign layer_1_weights[15][122] = 6'sd3;
    assign layer_1_weights[15][123] = 6'sd5;
    assign layer_1_weights[15][124] = 6'sd3;
    assign layer_1_weights[15][125] = 6'sd1;
    assign layer_1_weights[15][126] = 6'sd0;
    assign layer_1_weights[15][127] = 6'sd3;
    assign layer_1_weights[15][128] = 6'sd2;
    assign layer_1_weights[15][129] = 6'sd3;
    assign layer_1_weights[15][130] = 6'sd2;
    assign layer_1_weights[15][131] = 6'sd8;
    assign layer_1_weights[15][132] = -6'sd1;
    assign layer_1_weights[15][133] = 6'sd10;
    assign layer_1_weights[15][134] = -6'sd8;
    assign layer_1_weights[15][135] = 6'sd0;
    assign layer_1_weights[15][136] = 6'sd3;
    assign layer_1_weights[15][137] = -6'sd3;
    assign layer_1_weights[15][138] = 6'sd2;
    assign layer_1_weights[15][139] = 6'sd3;
    assign layer_1_weights[15][140] = -6'sd1;
    assign layer_1_weights[15][141] = -6'sd7;
    assign layer_1_weights[15][142] = -6'sd1;
    assign layer_1_weights[15][143] = 6'sd1;
    assign layer_1_biases[15] = -6'sd4;
    assign layer_1_weights[16][0] = -6'sd1;
    assign layer_1_weights[16][1] = -6'sd1;
    assign layer_1_weights[16][2] = 6'sd3;
    assign layer_1_weights[16][3] = 6'sd11;
    assign layer_1_weights[16][4] = 6'sd18;
    assign layer_1_weights[16][5] = 6'sd12;
    assign layer_1_weights[16][6] = -6'sd1;
    assign layer_1_weights[16][7] = 6'sd4;
    assign layer_1_weights[16][8] = 6'sd11;
    assign layer_1_weights[16][9] = 6'sd12;
    assign layer_1_weights[16][10] = -6'sd1;
    assign layer_1_weights[16][11] = 6'sd0;
    assign layer_1_weights[16][12] = 6'sd1;
    assign layer_1_weights[16][13] = 6'sd0;
    assign layer_1_weights[16][14] = 6'sd3;
    assign layer_1_weights[16][15] = 6'sd5;
    assign layer_1_weights[16][16] = 6'sd9;
    assign layer_1_weights[16][17] = 6'sd3;
    assign layer_1_weights[16][18] = -6'sd1;
    assign layer_1_weights[16][19] = 6'sd2;
    assign layer_1_weights[16][20] = 6'sd5;
    assign layer_1_weights[16][21] = 6'sd8;
    assign layer_1_weights[16][22] = 6'sd2;
    assign layer_1_weights[16][23] = 6'sd0;
    assign layer_1_weights[16][24] = 6'sd2;
    assign layer_1_weights[16][25] = 6'sd1;
    assign layer_1_weights[16][26] = 6'sd9;
    assign layer_1_weights[16][27] = 6'sd2;
    assign layer_1_weights[16][28] = 6'sd3;
    assign layer_1_weights[16][29] = -6'sd2;
    assign layer_1_weights[16][30] = -6'sd3;
    assign layer_1_weights[16][31] = 6'sd1;
    assign layer_1_weights[16][32] = 6'sd2;
    assign layer_1_weights[16][33] = -6'sd2;
    assign layer_1_weights[16][34] = 6'sd5;
    assign layer_1_weights[16][35] = 6'sd6;
    assign layer_1_weights[16][36] = 6'sd2;
    assign layer_1_weights[16][37] = 6'sd2;
    assign layer_1_weights[16][38] = 6'sd0;
    assign layer_1_weights[16][39] = 6'sd2;
    assign layer_1_weights[16][40] = 6'sd7;
    assign layer_1_weights[16][41] = 6'sd1;
    assign layer_1_weights[16][42] = -6'sd2;
    assign layer_1_weights[16][43] = -6'sd2;
    assign layer_1_weights[16][44] = -6'sd1;
    assign layer_1_weights[16][45] = -6'sd4;
    assign layer_1_weights[16][46] = 6'sd0;
    assign layer_1_weights[16][47] = 6'sd5;
    assign layer_1_weights[16][48] = 6'sd2;
    assign layer_1_weights[16][49] = -6'sd2;
    assign layer_1_weights[16][50] = 6'sd0;
    assign layer_1_weights[16][51] = 6'sd3;
    assign layer_1_weights[16][52] = -6'sd1;
    assign layer_1_weights[16][53] = -6'sd2;
    assign layer_1_weights[16][54] = 6'sd0;
    assign layer_1_weights[16][55] = -6'sd2;
    assign layer_1_weights[16][56] = -6'sd5;
    assign layer_1_weights[16][57] = -6'sd2;
    assign layer_1_weights[16][58] = -6'sd4;
    assign layer_1_weights[16][59] = 6'sd3;
    assign layer_1_weights[16][60] = 6'sd2;
    assign layer_1_weights[16][61] = -6'sd9;
    assign layer_1_weights[16][62] = -6'sd8;
    assign layer_1_weights[16][63] = -6'sd5;
    assign layer_1_weights[16][64] = -6'sd9;
    assign layer_1_weights[16][65] = -6'sd5;
    assign layer_1_weights[16][66] = 6'sd2;
    assign layer_1_weights[16][67] = -6'sd2;
    assign layer_1_weights[16][68] = 6'sd1;
    assign layer_1_weights[16][69] = 6'sd1;
    assign layer_1_weights[16][70] = 6'sd6;
    assign layer_1_weights[16][71] = 6'sd4;
    assign layer_1_weights[16][72] = -6'sd6;
    assign layer_1_weights[16][73] = -6'sd8;
    assign layer_1_weights[16][74] = -6'sd5;
    assign layer_1_weights[16][75] = -6'sd8;
    assign layer_1_weights[16][76] = -6'sd3;
    assign layer_1_weights[16][77] = 6'sd7;
    assign layer_1_weights[16][78] = 6'sd4;
    assign layer_1_weights[16][79] = -6'sd3;
    assign layer_1_weights[16][80] = 6'sd3;
    assign layer_1_weights[16][81] = 6'sd3;
    assign layer_1_weights[16][82] = -6'sd1;
    assign layer_1_weights[16][83] = 6'sd7;
    assign layer_1_weights[16][84] = -6'sd7;
    assign layer_1_weights[16][85] = -6'sd6;
    assign layer_1_weights[16][86] = 6'sd1;
    assign layer_1_weights[16][87] = -6'sd1;
    assign layer_1_weights[16][88] = 6'sd3;
    assign layer_1_weights[16][89] = 6'sd8;
    assign layer_1_weights[16][90] = 6'sd2;
    assign layer_1_weights[16][91] = -6'sd1;
    assign layer_1_weights[16][92] = 6'sd0;
    assign layer_1_weights[16][93] = 6'sd0;
    assign layer_1_weights[16][94] = 6'sd2;
    assign layer_1_weights[16][95] = 6'sd3;
    assign layer_1_weights[16][96] = -6'sd3;
    assign layer_1_weights[16][97] = -6'sd1;
    assign layer_1_weights[16][98] = 6'sd3;
    assign layer_1_weights[16][99] = 6'sd1;
    assign layer_1_weights[16][100] = 6'sd4;
    assign layer_1_weights[16][101] = 6'sd4;
    assign layer_1_weights[16][102] = 6'sd0;
    assign layer_1_weights[16][103] = 6'sd3;
    assign layer_1_weights[16][104] = -6'sd1;
    assign layer_1_weights[16][105] = -6'sd1;
    assign layer_1_weights[16][106] = 6'sd0;
    assign layer_1_weights[16][107] = 6'sd13;
    assign layer_1_weights[16][108] = 6'sd9;
    assign layer_1_weights[16][109] = 6'sd2;
    assign layer_1_weights[16][110] = -6'sd3;
    assign layer_1_weights[16][111] = -6'sd1;
    assign layer_1_weights[16][112] = 6'sd4;
    assign layer_1_weights[16][113] = 6'sd5;
    assign layer_1_weights[16][114] = 6'sd4;
    assign layer_1_weights[16][115] = 6'sd1;
    assign layer_1_weights[16][116] = -6'sd2;
    assign layer_1_weights[16][117] = 6'sd0;
    assign layer_1_weights[16][118] = -6'sd8;
    assign layer_1_weights[16][119] = 6'sd3;
    assign layer_1_weights[16][120] = 6'sd0;
    assign layer_1_weights[16][121] = 6'sd2;
    assign layer_1_weights[16][122] = 6'sd0;
    assign layer_1_weights[16][123] = -6'sd3;
    assign layer_1_weights[16][124] = -6'sd1;
    assign layer_1_weights[16][125] = -6'sd2;
    assign layer_1_weights[16][126] = 6'sd0;
    assign layer_1_weights[16][127] = -6'sd4;
    assign layer_1_weights[16][128] = -6'sd2;
    assign layer_1_weights[16][129] = -6'sd7;
    assign layer_1_weights[16][130] = -6'sd3;
    assign layer_1_weights[16][131] = 6'sd7;
    assign layer_1_weights[16][132] = 6'sd2;
    assign layer_1_weights[16][133] = 6'sd2;
    assign layer_1_weights[16][134] = -6'sd2;
    assign layer_1_weights[16][135] = -6'sd1;
    assign layer_1_weights[16][136] = 6'sd0;
    assign layer_1_weights[16][137] = -6'sd2;
    assign layer_1_weights[16][138] = -6'sd1;
    assign layer_1_weights[16][139] = -6'sd3;
    assign layer_1_weights[16][140] = -6'sd3;
    assign layer_1_weights[16][141] = -6'sd1;
    assign layer_1_weights[16][142] = 6'sd0;
    assign layer_1_weights[16][143] = -6'sd1;
    assign layer_1_biases[16] = 6'sd1;
    assign layer_1_weights[17][0] = 6'sd0;
    assign layer_1_weights[17][1] = -6'sd1;
    assign layer_1_weights[17][2] = -6'sd3;
    assign layer_1_weights[17][3] = -6'sd7;
    assign layer_1_weights[17][4] = -6'sd11;
    assign layer_1_weights[17][5] = -6'sd1;
    assign layer_1_weights[17][6] = -6'sd4;
    assign layer_1_weights[17][7] = 6'sd6;
    assign layer_1_weights[17][8] = -6'sd17;
    assign layer_1_weights[17][9] = -6'sd8;
    assign layer_1_weights[17][10] = 6'sd1;
    assign layer_1_weights[17][11] = 6'sd2;
    assign layer_1_weights[17][12] = -6'sd1;
    assign layer_1_weights[17][13] = -6'sd2;
    assign layer_1_weights[17][14] = -6'sd10;
    assign layer_1_weights[17][15] = -6'sd3;
    assign layer_1_weights[17][16] = -6'sd6;
    assign layer_1_weights[17][17] = -6'sd2;
    assign layer_1_weights[17][18] = -6'sd1;
    assign layer_1_weights[17][19] = -6'sd3;
    assign layer_1_weights[17][20] = -6'sd9;
    assign layer_1_weights[17][21] = -6'sd6;
    assign layer_1_weights[17][22] = -6'sd1;
    assign layer_1_weights[17][23] = -6'sd2;
    assign layer_1_weights[17][24] = 6'sd1;
    assign layer_1_weights[17][25] = -6'sd6;
    assign layer_1_weights[17][26] = -6'sd1;
    assign layer_1_weights[17][27] = -6'sd8;
    assign layer_1_weights[17][28] = -6'sd6;
    assign layer_1_weights[17][29] = -6'sd7;
    assign layer_1_weights[17][30] = -6'sd9;
    assign layer_1_weights[17][31] = -6'sd2;
    assign layer_1_weights[17][32] = 6'sd3;
    assign layer_1_weights[17][33] = -6'sd2;
    assign layer_1_weights[17][34] = 6'sd0;
    assign layer_1_weights[17][35] = -6'sd3;
    assign layer_1_weights[17][36] = 6'sd1;
    assign layer_1_weights[17][37] = -6'sd8;
    assign layer_1_weights[17][38] = 6'sd3;
    assign layer_1_weights[17][39] = 6'sd3;
    assign layer_1_weights[17][40] = 6'sd3;
    assign layer_1_weights[17][41] = -6'sd2;
    assign layer_1_weights[17][42] = 6'sd3;
    assign layer_1_weights[17][43] = 6'sd1;
    assign layer_1_weights[17][44] = 6'sd1;
    assign layer_1_weights[17][45] = 6'sd4;
    assign layer_1_weights[17][46] = 6'sd2;
    assign layer_1_weights[17][47] = -6'sd5;
    assign layer_1_weights[17][48] = -6'sd8;
    assign layer_1_weights[17][49] = -6'sd2;
    assign layer_1_weights[17][50] = 6'sd3;
    assign layer_1_weights[17][51] = 6'sd1;
    assign layer_1_weights[17][52] = 6'sd4;
    assign layer_1_weights[17][53] = 6'sd2;
    assign layer_1_weights[17][54] = 6'sd2;
    assign layer_1_weights[17][55] = 6'sd0;
    assign layer_1_weights[17][56] = -6'sd4;
    assign layer_1_weights[17][57] = 6'sd3;
    assign layer_1_weights[17][58] = 6'sd0;
    assign layer_1_weights[17][59] = -6'sd1;
    assign layer_1_weights[17][60] = -6'sd1;
    assign layer_1_weights[17][61] = 6'sd4;
    assign layer_1_weights[17][62] = 6'sd0;
    assign layer_1_weights[17][63] = -6'sd2;
    assign layer_1_weights[17][64] = 6'sd2;
    assign layer_1_weights[17][65] = 6'sd4;
    assign layer_1_weights[17][66] = -6'sd3;
    assign layer_1_weights[17][67] = -6'sd2;
    assign layer_1_weights[17][68] = -6'sd2;
    assign layer_1_weights[17][69] = 6'sd1;
    assign layer_1_weights[17][70] = 6'sd5;
    assign layer_1_weights[17][71] = 6'sd3;
    assign layer_1_weights[17][72] = -6'sd1;
    assign layer_1_weights[17][73] = -6'sd5;
    assign layer_1_weights[17][74] = -6'sd3;
    assign layer_1_weights[17][75] = -6'sd1;
    assign layer_1_weights[17][76] = 6'sd1;
    assign layer_1_weights[17][77] = 6'sd2;
    assign layer_1_weights[17][78] = 6'sd1;
    assign layer_1_weights[17][79] = 6'sd5;
    assign layer_1_weights[17][80] = 6'sd4;
    assign layer_1_weights[17][81] = 6'sd0;
    assign layer_1_weights[17][82] = 6'sd5;
    assign layer_1_weights[17][83] = 6'sd3;
    assign layer_1_weights[17][84] = -6'sd2;
    assign layer_1_weights[17][85] = 6'sd0;
    assign layer_1_weights[17][86] = 6'sd0;
    assign layer_1_weights[17][87] = 6'sd0;
    assign layer_1_weights[17][88] = 6'sd1;
    assign layer_1_weights[17][89] = 6'sd0;
    assign layer_1_weights[17][90] = 6'sd5;
    assign layer_1_weights[17][91] = 6'sd4;
    assign layer_1_weights[17][92] = 6'sd2;
    assign layer_1_weights[17][93] = 6'sd2;
    assign layer_1_weights[17][94] = 6'sd1;
    assign layer_1_weights[17][95] = 6'sd0;
    assign layer_1_weights[17][96] = 6'sd6;
    assign layer_1_weights[17][97] = -6'sd1;
    assign layer_1_weights[17][98] = -6'sd2;
    assign layer_1_weights[17][99] = 6'sd5;
    assign layer_1_weights[17][100] = 6'sd1;
    assign layer_1_weights[17][101] = 6'sd0;
    assign layer_1_weights[17][102] = -6'sd1;
    assign layer_1_weights[17][103] = -6'sd5;
    assign layer_1_weights[17][104] = 6'sd0;
    assign layer_1_weights[17][105] = -6'sd1;
    assign layer_1_weights[17][106] = -6'sd2;
    assign layer_1_weights[17][107] = 6'sd12;
    assign layer_1_weights[17][108] = -6'sd2;
    assign layer_1_weights[17][109] = 6'sd5;
    assign layer_1_weights[17][110] = 6'sd1;
    assign layer_1_weights[17][111] = -6'sd5;
    assign layer_1_weights[17][112] = -6'sd1;
    assign layer_1_weights[17][113] = -6'sd5;
    assign layer_1_weights[17][114] = -6'sd10;
    assign layer_1_weights[17][115] = -6'sd12;
    assign layer_1_weights[17][116] = -6'sd11;
    assign layer_1_weights[17][117] = -6'sd12;
    assign layer_1_weights[17][118] = -6'sd10;
    assign layer_1_weights[17][119] = 6'sd3;
    assign layer_1_weights[17][120] = 6'sd2;
    assign layer_1_weights[17][121] = -6'sd2;
    assign layer_1_weights[17][122] = -6'sd14;
    assign layer_1_weights[17][123] = -6'sd12;
    assign layer_1_weights[17][124] = -6'sd12;
    assign layer_1_weights[17][125] = -6'sd16;
    assign layer_1_weights[17][126] = -6'sd5;
    assign layer_1_weights[17][127] = 6'sd0;
    assign layer_1_weights[17][128] = -6'sd12;
    assign layer_1_weights[17][129] = -6'sd10;
    assign layer_1_weights[17][130] = -6'sd2;
    assign layer_1_weights[17][131] = 6'sd2;
    assign layer_1_weights[17][132] = -6'sd1;
    assign layer_1_weights[17][133] = 6'sd2;
    assign layer_1_weights[17][134] = -6'sd9;
    assign layer_1_weights[17][135] = -6'sd12;
    assign layer_1_weights[17][136] = -6'sd8;
    assign layer_1_weights[17][137] = 6'sd0;
    assign layer_1_weights[17][138] = -6'sd7;
    assign layer_1_weights[17][139] = -6'sd11;
    assign layer_1_weights[17][140] = 6'sd2;
    assign layer_1_weights[17][141] = 6'sd9;
    assign layer_1_weights[17][142] = 6'sd1;
    assign layer_1_weights[17][143] = 6'sd0;
    assign layer_1_biases[17] = 6'sd3;
    assign layer_1_weights[18][0] = 6'sd0;
    assign layer_1_weights[18][1] = -6'sd1;
    assign layer_1_weights[18][2] = 6'sd0;
    assign layer_1_weights[18][3] = 6'sd2;
    assign layer_1_weights[18][4] = 6'sd4;
    assign layer_1_weights[18][5] = 6'sd6;
    assign layer_1_weights[18][6] = -6'sd5;
    assign layer_1_weights[18][7] = -6'sd8;
    assign layer_1_weights[18][8] = 6'sd4;
    assign layer_1_weights[18][9] = -6'sd1;
    assign layer_1_weights[18][10] = 6'sd0;
    assign layer_1_weights[18][11] = 6'sd0;
    assign layer_1_weights[18][12] = 6'sd1;
    assign layer_1_weights[18][13] = 6'sd1;
    assign layer_1_weights[18][14] = -6'sd1;
    assign layer_1_weights[18][15] = -6'sd3;
    assign layer_1_weights[18][16] = 6'sd2;
    assign layer_1_weights[18][17] = -6'sd1;
    assign layer_1_weights[18][18] = 6'sd0;
    assign layer_1_weights[18][19] = 6'sd2;
    assign layer_1_weights[18][20] = 6'sd1;
    assign layer_1_weights[18][21] = 6'sd2;
    assign layer_1_weights[18][22] = 6'sd2;
    assign layer_1_weights[18][23] = -6'sd1;
    assign layer_1_weights[18][24] = -6'sd1;
    assign layer_1_weights[18][25] = 6'sd3;
    assign layer_1_weights[18][26] = -6'sd4;
    assign layer_1_weights[18][27] = -6'sd5;
    assign layer_1_weights[18][28] = 6'sd1;
    assign layer_1_weights[18][29] = 6'sd1;
    assign layer_1_weights[18][30] = -6'sd1;
    assign layer_1_weights[18][31] = 6'sd5;
    assign layer_1_weights[18][32] = 6'sd3;
    assign layer_1_weights[18][33] = -6'sd1;
    assign layer_1_weights[18][34] = -6'sd3;
    assign layer_1_weights[18][35] = -6'sd14;
    assign layer_1_weights[18][36] = -6'sd2;
    assign layer_1_weights[18][37] = 6'sd4;
    assign layer_1_weights[18][38] = 6'sd0;
    assign layer_1_weights[18][39] = 6'sd0;
    assign layer_1_weights[18][40] = 6'sd2;
    assign layer_1_weights[18][41] = -6'sd4;
    assign layer_1_weights[18][42] = -6'sd3;
    assign layer_1_weights[18][43] = 6'sd1;
    assign layer_1_weights[18][44] = 6'sd7;
    assign layer_1_weights[18][45] = -6'sd1;
    assign layer_1_weights[18][46] = 6'sd1;
    assign layer_1_weights[18][47] = -6'sd11;
    assign layer_1_weights[18][48] = -6'sd4;
    assign layer_1_weights[18][49] = 6'sd6;
    assign layer_1_weights[18][50] = -6'sd1;
    assign layer_1_weights[18][51] = 6'sd0;
    assign layer_1_weights[18][52] = -6'sd2;
    assign layer_1_weights[18][53] = -6'sd3;
    assign layer_1_weights[18][54] = -6'sd2;
    assign layer_1_weights[18][55] = -6'sd3;
    assign layer_1_weights[18][56] = -6'sd1;
    assign layer_1_weights[18][57] = 6'sd6;
    assign layer_1_weights[18][58] = 6'sd7;
    assign layer_1_weights[18][59] = 6'sd1;
    assign layer_1_weights[18][60] = -6'sd4;
    assign layer_1_weights[18][61] = -6'sd1;
    assign layer_1_weights[18][62] = 6'sd1;
    assign layer_1_weights[18][63] = 6'sd3;
    assign layer_1_weights[18][64] = 6'sd2;
    assign layer_1_weights[18][65] = -6'sd1;
    assign layer_1_weights[18][66] = -6'sd3;
    assign layer_1_weights[18][67] = -6'sd11;
    assign layer_1_weights[18][68] = -6'sd3;
    assign layer_1_weights[18][69] = 6'sd5;
    assign layer_1_weights[18][70] = 6'sd4;
    assign layer_1_weights[18][71] = 6'sd3;
    assign layer_1_weights[18][72] = 6'sd1;
    assign layer_1_weights[18][73] = 6'sd0;
    assign layer_1_weights[18][74] = 6'sd2;
    assign layer_1_weights[18][75] = 6'sd7;
    assign layer_1_weights[18][76] = 6'sd1;
    assign layer_1_weights[18][77] = -6'sd3;
    assign layer_1_weights[18][78] = -6'sd1;
    assign layer_1_weights[18][79] = -6'sd2;
    assign layer_1_weights[18][80] = 6'sd4;
    assign layer_1_weights[18][81] = 6'sd5;
    assign layer_1_weights[18][82] = 6'sd2;
    assign layer_1_weights[18][83] = -6'sd4;
    assign layer_1_weights[18][84] = -6'sd1;
    assign layer_1_weights[18][85] = 6'sd4;
    assign layer_1_weights[18][86] = 6'sd6;
    assign layer_1_weights[18][87] = 6'sd6;
    assign layer_1_weights[18][88] = -6'sd4;
    assign layer_1_weights[18][89] = -6'sd4;
    assign layer_1_weights[18][90] = -6'sd2;
    assign layer_1_weights[18][91] = 6'sd2;
    assign layer_1_weights[18][92] = 6'sd3;
    assign layer_1_weights[18][93] = 6'sd2;
    assign layer_1_weights[18][94] = 6'sd2;
    assign layer_1_weights[18][95] = 6'sd1;
    assign layer_1_weights[18][96] = -6'sd1;
    assign layer_1_weights[18][97] = 6'sd2;
    assign layer_1_weights[18][98] = 6'sd6;
    assign layer_1_weights[18][99] = 6'sd8;
    assign layer_1_weights[18][100] = -6'sd6;
    assign layer_1_weights[18][101] = -6'sd4;
    assign layer_1_weights[18][102] = 6'sd0;
    assign layer_1_weights[18][103] = -6'sd1;
    assign layer_1_weights[18][104] = 6'sd2;
    assign layer_1_weights[18][105] = 6'sd2;
    assign layer_1_weights[18][106] = -6'sd3;
    assign layer_1_weights[18][107] = -6'sd5;
    assign layer_1_weights[18][108] = -6'sd1;
    assign layer_1_weights[18][109] = 6'sd5;
    assign layer_1_weights[18][110] = 6'sd5;
    assign layer_1_weights[18][111] = 6'sd3;
    assign layer_1_weights[18][112] = 6'sd4;
    assign layer_1_weights[18][113] = -6'sd2;
    assign layer_1_weights[18][114] = -6'sd2;
    assign layer_1_weights[18][115] = -6'sd2;
    assign layer_1_weights[18][116] = 6'sd0;
    assign layer_1_weights[18][117] = -6'sd1;
    assign layer_1_weights[18][118] = -6'sd1;
    assign layer_1_weights[18][119] = -6'sd4;
    assign layer_1_weights[18][120] = -6'sd1;
    assign layer_1_weights[18][121] = -6'sd6;
    assign layer_1_weights[18][122] = 6'sd3;
    assign layer_1_weights[18][123] = 6'sd5;
    assign layer_1_weights[18][124] = 6'sd3;
    assign layer_1_weights[18][125] = -6'sd2;
    assign layer_1_weights[18][126] = 6'sd0;
    assign layer_1_weights[18][127] = -6'sd2;
    assign layer_1_weights[18][128] = -6'sd5;
    assign layer_1_weights[18][129] = -6'sd4;
    assign layer_1_weights[18][130] = -6'sd5;
    assign layer_1_weights[18][131] = -6'sd1;
    assign layer_1_weights[18][132] = -6'sd1;
    assign layer_1_weights[18][133] = 6'sd0;
    assign layer_1_weights[18][134] = -6'sd1;
    assign layer_1_weights[18][135] = 6'sd4;
    assign layer_1_weights[18][136] = 6'sd2;
    assign layer_1_weights[18][137] = -6'sd6;
    assign layer_1_weights[18][138] = -6'sd14;
    assign layer_1_weights[18][139] = -6'sd9;
    assign layer_1_weights[18][140] = -6'sd1;
    assign layer_1_weights[18][141] = -6'sd3;
    assign layer_1_weights[18][142] = -6'sd1;
    assign layer_1_weights[18][143] = 6'sd0;
    assign layer_1_biases[18] = -6'sd3;
    assign layer_1_weights[19][0] = -6'sd1;
    assign layer_1_weights[19][1] = -6'sd1;
    assign layer_1_weights[19][2] = 6'sd1;
    assign layer_1_weights[19][3] = 6'sd5;
    assign layer_1_weights[19][4] = -6'sd4;
    assign layer_1_weights[19][5] = 6'sd10;
    assign layer_1_weights[19][6] = 6'sd10;
    assign layer_1_weights[19][7] = 6'sd4;
    assign layer_1_weights[19][8] = 6'sd5;
    assign layer_1_weights[19][9] = 6'sd4;
    assign layer_1_weights[19][10] = 6'sd0;
    assign layer_1_weights[19][11] = 6'sd0;
    assign layer_1_weights[19][12] = 6'sd1;
    assign layer_1_weights[19][13] = 6'sd0;
    assign layer_1_weights[19][14] = -6'sd3;
    assign layer_1_weights[19][15] = 6'sd1;
    assign layer_1_weights[19][16] = 6'sd0;
    assign layer_1_weights[19][17] = -6'sd4;
    assign layer_1_weights[19][18] = -6'sd5;
    assign layer_1_weights[19][19] = -6'sd5;
    assign layer_1_weights[19][20] = -6'sd13;
    assign layer_1_weights[19][21] = 6'sd2;
    assign layer_1_weights[19][22] = 6'sd3;
    assign layer_1_weights[19][23] = 6'sd5;
    assign layer_1_weights[19][24] = -6'sd1;
    assign layer_1_weights[19][25] = 6'sd3;
    assign layer_1_weights[19][26] = -6'sd5;
    assign layer_1_weights[19][27] = -6'sd1;
    assign layer_1_weights[19][28] = -6'sd5;
    assign layer_1_weights[19][29] = -6'sd7;
    assign layer_1_weights[19][30] = -6'sd4;
    assign layer_1_weights[19][31] = -6'sd1;
    assign layer_1_weights[19][32] = 6'sd0;
    assign layer_1_weights[19][33] = -6'sd3;
    assign layer_1_weights[19][34] = 6'sd0;
    assign layer_1_weights[19][35] = 6'sd4;
    assign layer_1_weights[19][36] = 6'sd7;
    assign layer_1_weights[19][37] = 6'sd1;
    assign layer_1_weights[19][38] = 6'sd3;
    assign layer_1_weights[19][39] = 6'sd1;
    assign layer_1_weights[19][40] = -6'sd3;
    assign layer_1_weights[19][41] = 6'sd5;
    assign layer_1_weights[19][42] = 6'sd5;
    assign layer_1_weights[19][43] = 6'sd1;
    assign layer_1_weights[19][44] = -6'sd2;
    assign layer_1_weights[19][45] = -6'sd2;
    assign layer_1_weights[19][46] = -6'sd7;
    assign layer_1_weights[19][47] = -6'sd7;
    assign layer_1_weights[19][48] = 6'sd12;
    assign layer_1_weights[19][49] = 6'sd5;
    assign layer_1_weights[19][50] = 6'sd2;
    assign layer_1_weights[19][51] = 6'sd5;
    assign layer_1_weights[19][52] = 6'sd6;
    assign layer_1_weights[19][53] = 6'sd8;
    assign layer_1_weights[19][54] = 6'sd4;
    assign layer_1_weights[19][55] = 6'sd4;
    assign layer_1_weights[19][56] = 6'sd5;
    assign layer_1_weights[19][57] = 6'sd1;
    assign layer_1_weights[19][58] = 6'sd3;
    assign layer_1_weights[19][59] = 6'sd0;
    assign layer_1_weights[19][60] = 6'sd8;
    assign layer_1_weights[19][61] = 6'sd2;
    assign layer_1_weights[19][62] = 6'sd0;
    assign layer_1_weights[19][63] = 6'sd0;
    assign layer_1_weights[19][64] = -6'sd2;
    assign layer_1_weights[19][65] = 6'sd0;
    assign layer_1_weights[19][66] = 6'sd0;
    assign layer_1_weights[19][67] = 6'sd0;
    assign layer_1_weights[19][68] = 6'sd2;
    assign layer_1_weights[19][69] = 6'sd3;
    assign layer_1_weights[19][70] = 6'sd2;
    assign layer_1_weights[19][71] = 6'sd0;
    assign layer_1_weights[19][72] = 6'sd1;
    assign layer_1_weights[19][73] = 6'sd1;
    assign layer_1_weights[19][74] = -6'sd4;
    assign layer_1_weights[19][75] = -6'sd2;
    assign layer_1_weights[19][76] = 6'sd2;
    assign layer_1_weights[19][77] = -6'sd2;
    assign layer_1_weights[19][78] = -6'sd5;
    assign layer_1_weights[19][79] = -6'sd6;
    assign layer_1_weights[19][80] = -6'sd1;
    assign layer_1_weights[19][81] = 6'sd6;
    assign layer_1_weights[19][82] = 6'sd4;
    assign layer_1_weights[19][83] = -6'sd11;
    assign layer_1_weights[19][84] = -6'sd2;
    assign layer_1_weights[19][85] = -6'sd3;
    assign layer_1_weights[19][86] = 6'sd2;
    assign layer_1_weights[19][87] = -6'sd1;
    assign layer_1_weights[19][88] = 6'sd0;
    assign layer_1_weights[19][89] = 6'sd0;
    assign layer_1_weights[19][90] = -6'sd4;
    assign layer_1_weights[19][91] = -6'sd2;
    assign layer_1_weights[19][92] = 6'sd1;
    assign layer_1_weights[19][93] = 6'sd4;
    assign layer_1_weights[19][94] = 6'sd1;
    assign layer_1_weights[19][95] = -6'sd5;
    assign layer_1_weights[19][96] = 6'sd2;
    assign layer_1_weights[19][97] = -6'sd2;
    assign layer_1_weights[19][98] = -6'sd1;
    assign layer_1_weights[19][99] = -6'sd3;
    assign layer_1_weights[19][100] = -6'sd3;
    assign layer_1_weights[19][101] = -6'sd2;
    assign layer_1_weights[19][102] = -6'sd1;
    assign layer_1_weights[19][103] = 6'sd3;
    assign layer_1_weights[19][104] = 6'sd2;
    assign layer_1_weights[19][105] = 6'sd4;
    assign layer_1_weights[19][106] = 6'sd3;
    assign layer_1_weights[19][107] = 6'sd3;
    assign layer_1_weights[19][108] = -6'sd4;
    assign layer_1_weights[19][109] = 6'sd1;
    assign layer_1_weights[19][110] = -6'sd2;
    assign layer_1_weights[19][111] = -6'sd1;
    assign layer_1_weights[19][112] = -6'sd4;
    assign layer_1_weights[19][113] = 6'sd0;
    assign layer_1_weights[19][114] = 6'sd1;
    assign layer_1_weights[19][115] = 6'sd1;
    assign layer_1_weights[19][116] = -6'sd1;
    assign layer_1_weights[19][117] = 6'sd3;
    assign layer_1_weights[19][118] = 6'sd0;
    assign layer_1_weights[19][119] = 6'sd5;
    assign layer_1_weights[19][120] = -6'sd2;
    assign layer_1_weights[19][121] = 6'sd5;
    assign layer_1_weights[19][122] = 6'sd1;
    assign layer_1_weights[19][123] = -6'sd1;
    assign layer_1_weights[19][124] = 6'sd3;
    assign layer_1_weights[19][125] = 6'sd5;
    assign layer_1_weights[19][126] = 6'sd2;
    assign layer_1_weights[19][127] = 6'sd2;
    assign layer_1_weights[19][128] = -6'sd2;
    assign layer_1_weights[19][129] = -6'sd2;
    assign layer_1_weights[19][130] = 6'sd2;
    assign layer_1_weights[19][131] = 6'sd2;
    assign layer_1_weights[19][132] = 6'sd0;
    assign layer_1_weights[19][133] = 6'sd6;
    assign layer_1_weights[19][134] = -6'sd3;
    assign layer_1_weights[19][135] = 6'sd6;
    assign layer_1_weights[19][136] = 6'sd7;
    assign layer_1_weights[19][137] = 6'sd9;
    assign layer_1_weights[19][138] = 6'sd5;
    assign layer_1_weights[19][139] = 6'sd4;
    assign layer_1_weights[19][140] = 6'sd14;
    assign layer_1_weights[19][141] = 6'sd2;
    assign layer_1_weights[19][142] = -6'sd1;
    assign layer_1_weights[19][143] = 6'sd0;
    assign layer_1_biases[19] = -6'sd2;
    assign layer_1_weights[20][0] = 6'sd0;
    assign layer_1_weights[20][1] = 6'sd2;
    assign layer_1_weights[20][2] = 6'sd3;
    assign layer_1_weights[20][3] = 6'sd11;
    assign layer_1_weights[20][4] = 6'sd12;
    assign layer_1_weights[20][5] = 6'sd13;
    assign layer_1_weights[20][6] = 6'sd3;
    assign layer_1_weights[20][7] = 6'sd3;
    assign layer_1_weights[20][8] = 6'sd6;
    assign layer_1_weights[20][9] = 6'sd8;
    assign layer_1_weights[20][10] = 6'sd1;
    assign layer_1_weights[20][11] = 6'sd0;
    assign layer_1_weights[20][12] = 6'sd1;
    assign layer_1_weights[20][13] = 6'sd0;
    assign layer_1_weights[20][14] = -6'sd5;
    assign layer_1_weights[20][15] = 6'sd4;
    assign layer_1_weights[20][16] = 6'sd2;
    assign layer_1_weights[20][17] = 6'sd4;
    assign layer_1_weights[20][18] = 6'sd0;
    assign layer_1_weights[20][19] = 6'sd0;
    assign layer_1_weights[20][20] = 6'sd1;
    assign layer_1_weights[20][21] = 6'sd0;
    assign layer_1_weights[20][22] = -6'sd3;
    assign layer_1_weights[20][23] = 6'sd3;
    assign layer_1_weights[20][24] = 6'sd0;
    assign layer_1_weights[20][25] = -6'sd8;
    assign layer_1_weights[20][26] = -6'sd14;
    assign layer_1_weights[20][27] = 6'sd0;
    assign layer_1_weights[20][28] = 6'sd1;
    assign layer_1_weights[20][29] = 6'sd5;
    assign layer_1_weights[20][30] = 6'sd5;
    assign layer_1_weights[20][31] = -6'sd2;
    assign layer_1_weights[20][32] = -6'sd3;
    assign layer_1_weights[20][33] = -6'sd3;
    assign layer_1_weights[20][34] = 6'sd1;
    assign layer_1_weights[20][35] = 6'sd6;
    assign layer_1_weights[20][36] = -6'sd7;
    assign layer_1_weights[20][37] = -6'sd4;
    assign layer_1_weights[20][38] = -6'sd4;
    assign layer_1_weights[20][39] = 6'sd3;
    assign layer_1_weights[20][40] = 6'sd6;
    assign layer_1_weights[20][41] = 6'sd1;
    assign layer_1_weights[20][42] = -6'sd2;
    assign layer_1_weights[20][43] = 6'sd1;
    assign layer_1_weights[20][44] = -6'sd2;
    assign layer_1_weights[20][45] = -6'sd4;
    assign layer_1_weights[20][46] = 6'sd2;
    assign layer_1_weights[20][47] = 6'sd1;
    assign layer_1_weights[20][48] = -6'sd8;
    assign layer_1_weights[20][49] = -6'sd4;
    assign layer_1_weights[20][50] = 6'sd1;
    assign layer_1_weights[20][51] = 6'sd9;
    assign layer_1_weights[20][52] = 6'sd3;
    assign layer_1_weights[20][53] = -6'sd7;
    assign layer_1_weights[20][54] = -6'sd1;
    assign layer_1_weights[20][55] = 6'sd3;
    assign layer_1_weights[20][56] = 6'sd2;
    assign layer_1_weights[20][57] = 6'sd0;
    assign layer_1_weights[20][58] = -6'sd1;
    assign layer_1_weights[20][59] = -6'sd5;
    assign layer_1_weights[20][60] = -6'sd10;
    assign layer_1_weights[20][61] = -6'sd2;
    assign layer_1_weights[20][62] = 6'sd3;
    assign layer_1_weights[20][63] = 6'sd5;
    assign layer_1_weights[20][64] = 6'sd3;
    assign layer_1_weights[20][65] = 6'sd0;
    assign layer_1_weights[20][66] = -6'sd1;
    assign layer_1_weights[20][67] = 6'sd1;
    assign layer_1_weights[20][68] = -6'sd1;
    assign layer_1_weights[20][69] = 6'sd1;
    assign layer_1_weights[20][70] = 6'sd6;
    assign layer_1_weights[20][71] = 6'sd0;
    assign layer_1_weights[20][72] = -6'sd6;
    assign layer_1_weights[20][73] = 6'sd0;
    assign layer_1_weights[20][74] = 6'sd2;
    assign layer_1_weights[20][75] = 6'sd0;
    assign layer_1_weights[20][76] = 6'sd1;
    assign layer_1_weights[20][77] = 6'sd2;
    assign layer_1_weights[20][78] = -6'sd2;
    assign layer_1_weights[20][79] = 6'sd1;
    assign layer_1_weights[20][80] = -6'sd3;
    assign layer_1_weights[20][81] = -6'sd2;
    assign layer_1_weights[20][82] = 6'sd2;
    assign layer_1_weights[20][83] = 6'sd12;
    assign layer_1_weights[20][84] = -6'sd3;
    assign layer_1_weights[20][85] = 6'sd0;
    assign layer_1_weights[20][86] = 6'sd1;
    assign layer_1_weights[20][87] = -6'sd2;
    assign layer_1_weights[20][88] = 6'sd4;
    assign layer_1_weights[20][89] = 6'sd4;
    assign layer_1_weights[20][90] = -6'sd2;
    assign layer_1_weights[20][91] = -6'sd1;
    assign layer_1_weights[20][92] = -6'sd2;
    assign layer_1_weights[20][93] = -6'sd1;
    assign layer_1_weights[20][94] = -6'sd1;
    assign layer_1_weights[20][95] = 6'sd1;
    assign layer_1_weights[20][96] = 6'sd6;
    assign layer_1_weights[20][97] = -6'sd3;
    assign layer_1_weights[20][98] = -6'sd2;
    assign layer_1_weights[20][99] = -6'sd2;
    assign layer_1_weights[20][100] = 6'sd3;
    assign layer_1_weights[20][101] = -6'sd2;
    assign layer_1_weights[20][102] = -6'sd2;
    assign layer_1_weights[20][103] = 6'sd0;
    assign layer_1_weights[20][104] = 6'sd1;
    assign layer_1_weights[20][105] = 6'sd5;
    assign layer_1_weights[20][106] = 6'sd5;
    assign layer_1_weights[20][107] = 6'sd4;
    assign layer_1_weights[20][108] = 6'sd4;
    assign layer_1_weights[20][109] = 6'sd2;
    assign layer_1_weights[20][110] = -6'sd2;
    assign layer_1_weights[20][111] = -6'sd1;
    assign layer_1_weights[20][112] = 6'sd0;
    assign layer_1_weights[20][113] = 6'sd2;
    assign layer_1_weights[20][114] = 6'sd1;
    assign layer_1_weights[20][115] = -6'sd4;
    assign layer_1_weights[20][116] = 6'sd0;
    assign layer_1_weights[20][117] = 6'sd4;
    assign layer_1_weights[20][118] = 6'sd8;
    assign layer_1_weights[20][119] = -6'sd3;
    assign layer_1_weights[20][120] = 6'sd2;
    assign layer_1_weights[20][121] = 6'sd4;
    assign layer_1_weights[20][122] = -6'sd5;
    assign layer_1_weights[20][123] = -6'sd3;
    assign layer_1_weights[20][124] = -6'sd2;
    assign layer_1_weights[20][125] = -6'sd2;
    assign layer_1_weights[20][126] = -6'sd2;
    assign layer_1_weights[20][127] = 6'sd3;
    assign layer_1_weights[20][128] = 6'sd4;
    assign layer_1_weights[20][129] = 6'sd7;
    assign layer_1_weights[20][130] = 6'sd3;
    assign layer_1_weights[20][131] = -6'sd1;
    assign layer_1_weights[20][132] = 6'sd1;
    assign layer_1_weights[20][133] = 6'sd0;
    assign layer_1_weights[20][134] = -6'sd4;
    assign layer_1_weights[20][135] = 6'sd1;
    assign layer_1_weights[20][136] = -6'sd3;
    assign layer_1_weights[20][137] = -6'sd1;
    assign layer_1_weights[20][138] = -6'sd2;
    assign layer_1_weights[20][139] = -6'sd1;
    assign layer_1_weights[20][140] = -6'sd2;
    assign layer_1_weights[20][141] = -6'sd2;
    assign layer_1_weights[20][142] = -6'sd2;
    assign layer_1_weights[20][143] = 6'sd1;
    assign layer_1_biases[20] = -6'sd5;
    assign layer_1_weights[21][0] = 6'sd1;
    assign layer_1_weights[21][1] = -6'sd2;
    assign layer_1_weights[21][2] = 6'sd3;
    assign layer_1_weights[21][3] = -6'sd1;
    assign layer_1_weights[21][4] = 6'sd4;
    assign layer_1_weights[21][5] = 6'sd14;
    assign layer_1_weights[21][6] = 6'sd0;
    assign layer_1_weights[21][7] = 6'sd4;
    assign layer_1_weights[21][8] = 6'sd3;
    assign layer_1_weights[21][9] = 6'sd3;
    assign layer_1_weights[21][10] = 6'sd2;
    assign layer_1_weights[21][11] = 6'sd1;
    assign layer_1_weights[21][12] = 6'sd1;
    assign layer_1_weights[21][13] = -6'sd1;
    assign layer_1_weights[21][14] = -6'sd2;
    assign layer_1_weights[21][15] = -6'sd1;
    assign layer_1_weights[21][16] = -6'sd1;
    assign layer_1_weights[21][17] = -6'sd2;
    assign layer_1_weights[21][18] = -6'sd4;
    assign layer_1_weights[21][19] = 6'sd1;
    assign layer_1_weights[21][20] = -6'sd2;
    assign layer_1_weights[21][21] = -6'sd2;
    assign layer_1_weights[21][22] = 6'sd1;
    assign layer_1_weights[21][23] = 6'sd7;
    assign layer_1_weights[21][24] = 6'sd0;
    assign layer_1_weights[21][25] = 6'sd0;
    assign layer_1_weights[21][26] = -6'sd2;
    assign layer_1_weights[21][27] = 6'sd0;
    assign layer_1_weights[21][28] = 6'sd0;
    assign layer_1_weights[21][29] = 6'sd4;
    assign layer_1_weights[21][30] = 6'sd3;
    assign layer_1_weights[21][31] = 6'sd2;
    assign layer_1_weights[21][32] = 6'sd4;
    assign layer_1_weights[21][33] = 6'sd3;
    assign layer_1_weights[21][34] = 6'sd4;
    assign layer_1_weights[21][35] = 6'sd7;
    assign layer_1_weights[21][36] = -6'sd2;
    assign layer_1_weights[21][37] = -6'sd1;
    assign layer_1_weights[21][38] = -6'sd1;
    assign layer_1_weights[21][39] = 6'sd1;
    assign layer_1_weights[21][40] = 6'sd4;
    assign layer_1_weights[21][41] = 6'sd4;
    assign layer_1_weights[21][42] = 6'sd4;
    assign layer_1_weights[21][43] = 6'sd2;
    assign layer_1_weights[21][44] = 6'sd2;
    assign layer_1_weights[21][45] = 6'sd5;
    assign layer_1_weights[21][46] = 6'sd5;
    assign layer_1_weights[21][47] = 6'sd8;
    assign layer_1_weights[21][48] = 6'sd1;
    assign layer_1_weights[21][49] = 6'sd0;
    assign layer_1_weights[21][50] = 6'sd2;
    assign layer_1_weights[21][51] = 6'sd2;
    assign layer_1_weights[21][52] = -6'sd3;
    assign layer_1_weights[21][53] = -6'sd2;
    assign layer_1_weights[21][54] = -6'sd5;
    assign layer_1_weights[21][55] = -6'sd9;
    assign layer_1_weights[21][56] = -6'sd12;
    assign layer_1_weights[21][57] = -6'sd12;
    assign layer_1_weights[21][58] = -6'sd7;
    assign layer_1_weights[21][59] = -6'sd4;
    assign layer_1_weights[21][60] = -6'sd4;
    assign layer_1_weights[21][61] = 6'sd2;
    assign layer_1_weights[21][62] = 6'sd0;
    assign layer_1_weights[21][63] = 6'sd2;
    assign layer_1_weights[21][64] = 6'sd1;
    assign layer_1_weights[21][65] = 6'sd4;
    assign layer_1_weights[21][66] = -6'sd2;
    assign layer_1_weights[21][67] = -6'sd6;
    assign layer_1_weights[21][68] = -6'sd5;
    assign layer_1_weights[21][69] = -6'sd9;
    assign layer_1_weights[21][70] = -6'sd10;
    assign layer_1_weights[21][71] = 6'sd0;
    assign layer_1_weights[21][72] = -6'sd3;
    assign layer_1_weights[21][73] = -6'sd4;
    assign layer_1_weights[21][74] = -6'sd2;
    assign layer_1_weights[21][75] = 6'sd3;
    assign layer_1_weights[21][76] = 6'sd2;
    assign layer_1_weights[21][77] = 6'sd2;
    assign layer_1_weights[21][78] = 6'sd2;
    assign layer_1_weights[21][79] = 6'sd2;
    assign layer_1_weights[21][80] = 6'sd0;
    assign layer_1_weights[21][81] = 6'sd0;
    assign layer_1_weights[21][82] = 6'sd3;
    assign layer_1_weights[21][83] = -6'sd2;
    assign layer_1_weights[21][84] = -6'sd4;
    assign layer_1_weights[21][85] = -6'sd4;
    assign layer_1_weights[21][86] = -6'sd2;
    assign layer_1_weights[21][87] = -6'sd1;
    assign layer_1_weights[21][88] = -6'sd4;
    assign layer_1_weights[21][89] = 6'sd0;
    assign layer_1_weights[21][90] = 6'sd0;
    assign layer_1_weights[21][91] = 6'sd1;
    assign layer_1_weights[21][92] = 6'sd3;
    assign layer_1_weights[21][93] = 6'sd3;
    assign layer_1_weights[21][94] = -6'sd2;
    assign layer_1_weights[21][95] = -6'sd4;
    assign layer_1_weights[21][96] = -6'sd2;
    assign layer_1_weights[21][97] = 6'sd3;
    assign layer_1_weights[21][98] = 6'sd3;
    assign layer_1_weights[21][99] = 6'sd0;
    assign layer_1_weights[21][100] = -6'sd7;
    assign layer_1_weights[21][101] = -6'sd4;
    assign layer_1_weights[21][102] = -6'sd1;
    assign layer_1_weights[21][103] = 6'sd1;
    assign layer_1_weights[21][104] = 6'sd4;
    assign layer_1_weights[21][105] = 6'sd6;
    assign layer_1_weights[21][106] = 6'sd1;
    assign layer_1_weights[21][107] = -6'sd3;
    assign layer_1_weights[21][108] = 6'sd1;
    assign layer_1_weights[21][109] = 6'sd7;
    assign layer_1_weights[21][110] = 6'sd3;
    assign layer_1_weights[21][111] = 6'sd2;
    assign layer_1_weights[21][112] = 6'sd4;
    assign layer_1_weights[21][113] = 6'sd1;
    assign layer_1_weights[21][114] = 6'sd2;
    assign layer_1_weights[21][115] = 6'sd2;
    assign layer_1_weights[21][116] = 6'sd5;
    assign layer_1_weights[21][117] = 6'sd1;
    assign layer_1_weights[21][118] = 6'sd3;
    assign layer_1_weights[21][119] = 6'sd8;
    assign layer_1_weights[21][120] = -6'sd2;
    assign layer_1_weights[21][121] = 6'sd8;
    assign layer_1_weights[21][122] = 6'sd10;
    assign layer_1_weights[21][123] = 6'sd6;
    assign layer_1_weights[21][124] = 6'sd6;
    assign layer_1_weights[21][125] = 6'sd2;
    assign layer_1_weights[21][126] = 6'sd4;
    assign layer_1_weights[21][127] = 6'sd1;
    assign layer_1_weights[21][128] = 6'sd2;
    assign layer_1_weights[21][129] = 6'sd3;
    assign layer_1_weights[21][130] = 6'sd9;
    assign layer_1_weights[21][131] = -6'sd2;
    assign layer_1_weights[21][132] = 6'sd0;
    assign layer_1_weights[21][133] = -6'sd1;
    assign layer_1_weights[21][134] = 6'sd3;
    assign layer_1_weights[21][135] = 6'sd7;
    assign layer_1_weights[21][136] = 6'sd2;
    assign layer_1_weights[21][137] = -6'sd2;
    assign layer_1_weights[21][138] = 6'sd3;
    assign layer_1_weights[21][139] = 6'sd5;
    assign layer_1_weights[21][140] = 6'sd4;
    assign layer_1_weights[21][141] = -6'sd1;
    assign layer_1_weights[21][142] = -6'sd2;
    assign layer_1_weights[21][143] = -6'sd1;
    assign layer_1_biases[21] = -6'sd4;
    assign layer_1_weights[22][0] = -6'sd2;
    assign layer_1_weights[22][1] = -6'sd1;
    assign layer_1_weights[22][2] = -6'sd3;
    assign layer_1_weights[22][3] = -6'sd6;
    assign layer_1_weights[22][4] = -6'sd5;
    assign layer_1_weights[22][5] = -6'sd10;
    assign layer_1_weights[22][6] = -6'sd2;
    assign layer_1_weights[22][7] = -6'sd4;
    assign layer_1_weights[22][8] = -6'sd11;
    assign layer_1_weights[22][9] = -6'sd6;
    assign layer_1_weights[22][10] = 6'sd1;
    assign layer_1_weights[22][11] = 6'sd0;
    assign layer_1_weights[22][12] = -6'sd1;
    assign layer_1_weights[22][13] = -6'sd1;
    assign layer_1_weights[22][14] = -6'sd2;
    assign layer_1_weights[22][15] = 6'sd0;
    assign layer_1_weights[22][16] = -6'sd3;
    assign layer_1_weights[22][17] = 6'sd1;
    assign layer_1_weights[22][18] = -6'sd2;
    assign layer_1_weights[22][19] = -6'sd3;
    assign layer_1_weights[22][20] = -6'sd1;
    assign layer_1_weights[22][21] = 6'sd1;
    assign layer_1_weights[22][22] = 6'sd5;
    assign layer_1_weights[22][23] = -6'sd1;
    assign layer_1_weights[22][24] = 6'sd1;
    assign layer_1_weights[22][25] = -6'sd1;
    assign layer_1_weights[22][26] = -6'sd6;
    assign layer_1_weights[22][27] = -6'sd1;
    assign layer_1_weights[22][28] = 6'sd0;
    assign layer_1_weights[22][29] = 6'sd2;
    assign layer_1_weights[22][30] = 6'sd4;
    assign layer_1_weights[22][31] = 6'sd1;
    assign layer_1_weights[22][32] = -6'sd2;
    assign layer_1_weights[22][33] = 6'sd0;
    assign layer_1_weights[22][34] = 6'sd1;
    assign layer_1_weights[22][35] = 6'sd2;
    assign layer_1_weights[22][36] = -6'sd3;
    assign layer_1_weights[22][37] = -6'sd6;
    assign layer_1_weights[22][38] = 6'sd1;
    assign layer_1_weights[22][39] = 6'sd0;
    assign layer_1_weights[22][40] = 6'sd3;
    assign layer_1_weights[22][41] = -6'sd1;
    assign layer_1_weights[22][42] = -6'sd4;
    assign layer_1_weights[22][43] = -6'sd3;
    assign layer_1_weights[22][44] = -6'sd1;
    assign layer_1_weights[22][45] = 6'sd3;
    assign layer_1_weights[22][46] = 6'sd0;
    assign layer_1_weights[22][47] = 6'sd5;
    assign layer_1_weights[22][48] = -6'sd5;
    assign layer_1_weights[22][49] = 6'sd1;
    assign layer_1_weights[22][50] = -6'sd1;
    assign layer_1_weights[22][51] = 6'sd2;
    assign layer_1_weights[22][52] = 6'sd3;
    assign layer_1_weights[22][53] = 6'sd0;
    assign layer_1_weights[22][54] = -6'sd3;
    assign layer_1_weights[22][55] = -6'sd4;
    assign layer_1_weights[22][56] = 6'sd1;
    assign layer_1_weights[22][57] = 6'sd3;
    assign layer_1_weights[22][58] = 6'sd0;
    assign layer_1_weights[22][59] = -6'sd1;
    assign layer_1_weights[22][60] = 6'sd1;
    assign layer_1_weights[22][61] = 6'sd5;
    assign layer_1_weights[22][62] = 6'sd3;
    assign layer_1_weights[22][63] = 6'sd2;
    assign layer_1_weights[22][64] = 6'sd2;
    assign layer_1_weights[22][65] = 6'sd2;
    assign layer_1_weights[22][66] = 6'sd3;
    assign layer_1_weights[22][67] = 6'sd1;
    assign layer_1_weights[22][68] = 6'sd3;
    assign layer_1_weights[22][69] = 6'sd2;
    assign layer_1_weights[22][70] = 6'sd1;
    assign layer_1_weights[22][71] = 6'sd1;
    assign layer_1_weights[22][72] = 6'sd0;
    assign layer_1_weights[22][73] = -6'sd4;
    assign layer_1_weights[22][74] = 6'sd2;
    assign layer_1_weights[22][75] = 6'sd4;
    assign layer_1_weights[22][76] = 6'sd1;
    assign layer_1_weights[22][77] = 6'sd3;
    assign layer_1_weights[22][78] = 6'sd9;
    assign layer_1_weights[22][79] = 6'sd7;
    assign layer_1_weights[22][80] = 6'sd4;
    assign layer_1_weights[22][81] = 6'sd0;
    assign layer_1_weights[22][82] = 6'sd0;
    assign layer_1_weights[22][83] = 6'sd2;
    assign layer_1_weights[22][84] = -6'sd2;
    assign layer_1_weights[22][85] = -6'sd5;
    assign layer_1_weights[22][86] = 6'sd5;
    assign layer_1_weights[22][87] = 6'sd4;
    assign layer_1_weights[22][88] = 6'sd6;
    assign layer_1_weights[22][89] = 6'sd1;
    assign layer_1_weights[22][90] = 6'sd5;
    assign layer_1_weights[22][91] = 6'sd6;
    assign layer_1_weights[22][92] = 6'sd2;
    assign layer_1_weights[22][93] = 6'sd2;
    assign layer_1_weights[22][94] = 6'sd0;
    assign layer_1_weights[22][95] = 6'sd3;
    assign layer_1_weights[22][96] = -6'sd9;
    assign layer_1_weights[22][97] = -6'sd1;
    assign layer_1_weights[22][98] = 6'sd1;
    assign layer_1_weights[22][99] = 6'sd2;
    assign layer_1_weights[22][100] = -6'sd4;
    assign layer_1_weights[22][101] = -6'sd6;
    assign layer_1_weights[22][102] = 6'sd0;
    assign layer_1_weights[22][103] = 6'sd1;
    assign layer_1_weights[22][104] = -6'sd1;
    assign layer_1_weights[22][105] = -6'sd2;
    assign layer_1_weights[22][106] = -6'sd3;
    assign layer_1_weights[22][107] = -6'sd1;
    assign layer_1_weights[22][108] = -6'sd4;
    assign layer_1_weights[22][109] = 6'sd0;
    assign layer_1_weights[22][110] = 6'sd1;
    assign layer_1_weights[22][111] = 6'sd1;
    assign layer_1_weights[22][112] = 6'sd0;
    assign layer_1_weights[22][113] = -6'sd4;
    assign layer_1_weights[22][114] = -6'sd4;
    assign layer_1_weights[22][115] = -6'sd2;
    assign layer_1_weights[22][116] = -6'sd1;
    assign layer_1_weights[22][117] = 6'sd1;
    assign layer_1_weights[22][118] = -6'sd3;
    assign layer_1_weights[22][119] = -6'sd1;
    assign layer_1_weights[22][120] = 6'sd1;
    assign layer_1_weights[22][121] = -6'sd7;
    assign layer_1_weights[22][122] = -6'sd1;
    assign layer_1_weights[22][123] = -6'sd3;
    assign layer_1_weights[22][124] = -6'sd3;
    assign layer_1_weights[22][125] = -6'sd3;
    assign layer_1_weights[22][126] = -6'sd2;
    assign layer_1_weights[22][127] = 6'sd1;
    assign layer_1_weights[22][128] = 6'sd4;
    assign layer_1_weights[22][129] = 6'sd6;
    assign layer_1_weights[22][130] = -6'sd1;
    assign layer_1_weights[22][131] = -6'sd7;
    assign layer_1_weights[22][132] = 6'sd0;
    assign layer_1_weights[22][133] = 6'sd2;
    assign layer_1_weights[22][134] = 6'sd0;
    assign layer_1_weights[22][135] = 6'sd2;
    assign layer_1_weights[22][136] = 6'sd0;
    assign layer_1_weights[22][137] = 6'sd0;
    assign layer_1_weights[22][138] = 6'sd3;
    assign layer_1_weights[22][139] = 6'sd1;
    assign layer_1_weights[22][140] = 6'sd0;
    assign layer_1_weights[22][141] = 6'sd6;
    assign layer_1_weights[22][142] = 6'sd1;
    assign layer_1_weights[22][143] = 6'sd1;
    assign layer_1_biases[22] = 6'sd6;
    assign layer_1_weights[23][0] = -6'sd1;
    assign layer_1_weights[23][1] = -6'sd1;
    assign layer_1_weights[23][2] = 6'sd0;
    assign layer_1_weights[23][3] = -6'sd2;
    assign layer_1_weights[23][4] = 6'sd7;
    assign layer_1_weights[23][5] = -6'sd3;
    assign layer_1_weights[23][6] = 6'sd4;
    assign layer_1_weights[23][7] = -6'sd7;
    assign layer_1_weights[23][8] = 6'sd13;
    assign layer_1_weights[23][9] = 6'sd7;
    assign layer_1_weights[23][10] = 6'sd2;
    assign layer_1_weights[23][11] = 6'sd1;
    assign layer_1_weights[23][12] = 6'sd0;
    assign layer_1_weights[23][13] = 6'sd2;
    assign layer_1_weights[23][14] = -6'sd6;
    assign layer_1_weights[23][15] = -6'sd10;
    assign layer_1_weights[23][16] = -6'sd7;
    assign layer_1_weights[23][17] = -6'sd3;
    assign layer_1_weights[23][18] = -6'sd3;
    assign layer_1_weights[23][19] = -6'sd6;
    assign layer_1_weights[23][20] = -6'sd2;
    assign layer_1_weights[23][21] = -6'sd3;
    assign layer_1_weights[23][22] = 6'sd5;
    assign layer_1_weights[23][23] = -6'sd1;
    assign layer_1_weights[23][24] = 6'sd0;
    assign layer_1_weights[23][25] = -6'sd7;
    assign layer_1_weights[23][26] = -6'sd1;
    assign layer_1_weights[23][27] = -6'sd9;
    assign layer_1_weights[23][28] = -6'sd4;
    assign layer_1_weights[23][29] = -6'sd2;
    assign layer_1_weights[23][30] = 6'sd1;
    assign layer_1_weights[23][31] = 6'sd2;
    assign layer_1_weights[23][32] = 6'sd4;
    assign layer_1_weights[23][33] = 6'sd1;
    assign layer_1_weights[23][34] = 6'sd3;
    assign layer_1_weights[23][35] = 6'sd2;
    assign layer_1_weights[23][36] = 6'sd1;
    assign layer_1_weights[23][37] = 6'sd0;
    assign layer_1_weights[23][38] = 6'sd0;
    assign layer_1_weights[23][39] = -6'sd8;
    assign layer_1_weights[23][40] = -6'sd1;
    assign layer_1_weights[23][41] = 6'sd8;
    assign layer_1_weights[23][42] = 6'sd4;
    assign layer_1_weights[23][43] = -6'sd2;
    assign layer_1_weights[23][44] = 6'sd2;
    assign layer_1_weights[23][45] = 6'sd3;
    assign layer_1_weights[23][46] = -6'sd1;
    assign layer_1_weights[23][47] = 6'sd5;
    assign layer_1_weights[23][48] = 6'sd7;
    assign layer_1_weights[23][49] = -6'sd3;
    assign layer_1_weights[23][50] = -6'sd6;
    assign layer_1_weights[23][51] = -6'sd10;
    assign layer_1_weights[23][52] = 6'sd2;
    assign layer_1_weights[23][53] = 6'sd8;
    assign layer_1_weights[23][54] = -6'sd3;
    assign layer_1_weights[23][55] = -6'sd5;
    assign layer_1_weights[23][56] = -6'sd7;
    assign layer_1_weights[23][57] = -6'sd6;
    assign layer_1_weights[23][58] = 6'sd1;
    assign layer_1_weights[23][59] = 6'sd2;
    assign layer_1_weights[23][60] = 6'sd0;
    assign layer_1_weights[23][61] = 6'sd4;
    assign layer_1_weights[23][62] = -6'sd9;
    assign layer_1_weights[23][63] = -6'sd4;
    assign layer_1_weights[23][64] = 6'sd0;
    assign layer_1_weights[23][65] = 6'sd3;
    assign layer_1_weights[23][66] = 6'sd4;
    assign layer_1_weights[23][67] = 6'sd1;
    assign layer_1_weights[23][68] = -6'sd3;
    assign layer_1_weights[23][69] = 6'sd0;
    assign layer_1_weights[23][70] = -6'sd3;
    assign layer_1_weights[23][71] = -6'sd3;
    assign layer_1_weights[23][72] = 6'sd0;
    assign layer_1_weights[23][73] = 6'sd1;
    assign layer_1_weights[23][74] = -6'sd1;
    assign layer_1_weights[23][75] = -6'sd2;
    assign layer_1_weights[23][76] = -6'sd3;
    assign layer_1_weights[23][77] = 6'sd2;
    assign layer_1_weights[23][78] = 6'sd6;
    assign layer_1_weights[23][79] = 6'sd0;
    assign layer_1_weights[23][80] = 6'sd0;
    assign layer_1_weights[23][81] = 6'sd4;
    assign layer_1_weights[23][82] = 6'sd4;
    assign layer_1_weights[23][83] = -6'sd6;
    assign layer_1_weights[23][84] = -6'sd1;
    assign layer_1_weights[23][85] = 6'sd3;
    assign layer_1_weights[23][86] = 6'sd1;
    assign layer_1_weights[23][87] = 6'sd0;
    assign layer_1_weights[23][88] = -6'sd1;
    assign layer_1_weights[23][89] = 6'sd4;
    assign layer_1_weights[23][90] = 6'sd3;
    assign layer_1_weights[23][91] = -6'sd1;
    assign layer_1_weights[23][92] = 6'sd0;
    assign layer_1_weights[23][93] = 6'sd3;
    assign layer_1_weights[23][94] = -6'sd2;
    assign layer_1_weights[23][95] = -6'sd2;
    assign layer_1_weights[23][96] = -6'sd8;
    assign layer_1_weights[23][97] = -6'sd11;
    assign layer_1_weights[23][98] = -6'sd5;
    assign layer_1_weights[23][99] = 6'sd0;
    assign layer_1_weights[23][100] = 6'sd0;
    assign layer_1_weights[23][101] = 6'sd3;
    assign layer_1_weights[23][102] = 6'sd1;
    assign layer_1_weights[23][103] = -6'sd5;
    assign layer_1_weights[23][104] = -6'sd2;
    assign layer_1_weights[23][105] = -6'sd4;
    assign layer_1_weights[23][106] = 6'sd0;
    assign layer_1_weights[23][107] = 6'sd4;
    assign layer_1_weights[23][108] = -6'sd6;
    assign layer_1_weights[23][109] = -6'sd4;
    assign layer_1_weights[23][110] = -6'sd4;
    assign layer_1_weights[23][111] = -6'sd5;
    assign layer_1_weights[23][112] = 6'sd0;
    assign layer_1_weights[23][113] = 6'sd2;
    assign layer_1_weights[23][114] = -6'sd1;
    assign layer_1_weights[23][115] = -6'sd1;
    assign layer_1_weights[23][116] = -6'sd1;
    assign layer_1_weights[23][117] = -6'sd8;
    assign layer_1_weights[23][118] = 6'sd2;
    assign layer_1_weights[23][119] = 6'sd8;
    assign layer_1_weights[23][120] = 6'sd0;
    assign layer_1_weights[23][121] = -6'sd8;
    assign layer_1_weights[23][122] = -6'sd2;
    assign layer_1_weights[23][123] = -6'sd3;
    assign layer_1_weights[23][124] = -6'sd4;
    assign layer_1_weights[23][125] = 6'sd0;
    assign layer_1_weights[23][126] = 6'sd1;
    assign layer_1_weights[23][127] = 6'sd1;
    assign layer_1_weights[23][128] = -6'sd3;
    assign layer_1_weights[23][129] = -6'sd5;
    assign layer_1_weights[23][130] = 6'sd7;
    assign layer_1_weights[23][131] = -6'sd7;
    assign layer_1_weights[23][132] = -6'sd1;
    assign layer_1_weights[23][133] = 6'sd3;
    assign layer_1_weights[23][134] = 6'sd4;
    assign layer_1_weights[23][135] = 6'sd3;
    assign layer_1_weights[23][136] = 6'sd0;
    assign layer_1_weights[23][137] = 6'sd2;
    assign layer_1_weights[23][138] = 6'sd3;
    assign layer_1_weights[23][139] = 6'sd0;
    assign layer_1_weights[23][140] = 6'sd3;
    assign layer_1_weights[23][141] = 6'sd8;
    assign layer_1_weights[23][142] = 6'sd0;
    assign layer_1_weights[23][143] = -6'sd1;
    assign layer_1_biases[23] = 6'sd5;
    assign layer_1_weights[24][0] = 6'sd1;
    assign layer_1_weights[24][1] = -6'sd1;
    assign layer_1_weights[24][2] = 6'sd0;
    assign layer_1_weights[24][3] = 6'sd5;
    assign layer_1_weights[24][4] = 6'sd10;
    assign layer_1_weights[24][5] = 6'sd4;
    assign layer_1_weights[24][6] = 6'sd2;
    assign layer_1_weights[24][7] = -6'sd1;
    assign layer_1_weights[24][8] = -6'sd4;
    assign layer_1_weights[24][9] = -6'sd1;
    assign layer_1_weights[24][10] = 6'sd1;
    assign layer_1_weights[24][11] = 6'sd0;
    assign layer_1_weights[24][12] = 6'sd1;
    assign layer_1_weights[24][13] = 6'sd0;
    assign layer_1_weights[24][14] = -6'sd7;
    assign layer_1_weights[24][15] = -6'sd1;
    assign layer_1_weights[24][16] = -6'sd11;
    assign layer_1_weights[24][17] = -6'sd1;
    assign layer_1_weights[24][18] = -6'sd1;
    assign layer_1_weights[24][19] = -6'sd2;
    assign layer_1_weights[24][20] = 6'sd3;
    assign layer_1_weights[24][21] = 6'sd2;
    assign layer_1_weights[24][22] = 6'sd5;
    assign layer_1_weights[24][23] = 6'sd0;
    assign layer_1_weights[24][24] = -6'sd1;
    assign layer_1_weights[24][25] = 6'sd1;
    assign layer_1_weights[24][26] = -6'sd3;
    assign layer_1_weights[24][27] = -6'sd12;
    assign layer_1_weights[24][28] = 6'sd1;
    assign layer_1_weights[24][29] = 6'sd2;
    assign layer_1_weights[24][30] = 6'sd0;
    assign layer_1_weights[24][31] = -6'sd5;
    assign layer_1_weights[24][32] = -6'sd1;
    assign layer_1_weights[24][33] = 6'sd3;
    assign layer_1_weights[24][34] = 6'sd5;
    assign layer_1_weights[24][35] = 6'sd4;
    assign layer_1_weights[24][36] = -6'sd3;
    assign layer_1_weights[24][37] = -6'sd4;
    assign layer_1_weights[24][38] = -6'sd9;
    assign layer_1_weights[24][39] = -6'sd9;
    assign layer_1_weights[24][40] = -6'sd1;
    assign layer_1_weights[24][41] = 6'sd6;
    assign layer_1_weights[24][42] = -6'sd3;
    assign layer_1_weights[24][43] = 6'sd0;
    assign layer_1_weights[24][44] = 6'sd1;
    assign layer_1_weights[24][45] = 6'sd2;
    assign layer_1_weights[24][46] = 6'sd8;
    assign layer_1_weights[24][47] = 6'sd6;
    assign layer_1_weights[24][48] = -6'sd6;
    assign layer_1_weights[24][49] = 6'sd0;
    assign layer_1_weights[24][50] = -6'sd7;
    assign layer_1_weights[24][51] = -6'sd3;
    assign layer_1_weights[24][52] = 6'sd1;
    assign layer_1_weights[24][53] = 6'sd5;
    assign layer_1_weights[24][54] = -6'sd6;
    assign layer_1_weights[24][55] = -6'sd2;
    assign layer_1_weights[24][56] = 6'sd0;
    assign layer_1_weights[24][57] = -6'sd3;
    assign layer_1_weights[24][58] = 6'sd1;
    assign layer_1_weights[24][59] = 6'sd1;
    assign layer_1_weights[24][60] = 6'sd0;
    assign layer_1_weights[24][61] = -6'sd10;
    assign layer_1_weights[24][62] = -6'sd1;
    assign layer_1_weights[24][63] = -6'sd3;
    assign layer_1_weights[24][64] = 6'sd4;
    assign layer_1_weights[24][65] = 6'sd4;
    assign layer_1_weights[24][66] = -6'sd4;
    assign layer_1_weights[24][67] = -6'sd1;
    assign layer_1_weights[24][68] = -6'sd1;
    assign layer_1_weights[24][69] = -6'sd1;
    assign layer_1_weights[24][70] = 6'sd3;
    assign layer_1_weights[24][71] = -6'sd2;
    assign layer_1_weights[24][72] = -6'sd2;
    assign layer_1_weights[24][73] = -6'sd5;
    assign layer_1_weights[24][74] = -6'sd4;
    assign layer_1_weights[24][75] = 6'sd2;
    assign layer_1_weights[24][76] = 6'sd4;
    assign layer_1_weights[24][77] = 6'sd6;
    assign layer_1_weights[24][78] = -6'sd5;
    assign layer_1_weights[24][79] = 6'sd2;
    assign layer_1_weights[24][80] = 6'sd3;
    assign layer_1_weights[24][81] = 6'sd4;
    assign layer_1_weights[24][82] = 6'sd5;
    assign layer_1_weights[24][83] = -6'sd11;
    assign layer_1_weights[24][84] = -6'sd4;
    assign layer_1_weights[24][85] = -6'sd5;
    assign layer_1_weights[24][86] = 6'sd0;
    assign layer_1_weights[24][87] = 6'sd3;
    assign layer_1_weights[24][88] = 6'sd6;
    assign layer_1_weights[24][89] = -6'sd1;
    assign layer_1_weights[24][90] = 6'sd3;
    assign layer_1_weights[24][91] = 6'sd2;
    assign layer_1_weights[24][92] = -6'sd2;
    assign layer_1_weights[24][93] = 6'sd4;
    assign layer_1_weights[24][94] = -6'sd1;
    assign layer_1_weights[24][95] = -6'sd4;
    assign layer_1_weights[24][96] = 6'sd4;
    assign layer_1_weights[24][97] = 6'sd2;
    assign layer_1_weights[24][98] = -6'sd1;
    assign layer_1_weights[24][99] = 6'sd4;
    assign layer_1_weights[24][100] = 6'sd3;
    assign layer_1_weights[24][101] = -6'sd5;
    assign layer_1_weights[24][102] = -6'sd1;
    assign layer_1_weights[24][103] = -6'sd2;
    assign layer_1_weights[24][104] = -6'sd2;
    assign layer_1_weights[24][105] = -6'sd4;
    assign layer_1_weights[24][106] = -6'sd4;
    assign layer_1_weights[24][107] = -6'sd6;
    assign layer_1_weights[24][108] = -6'sd1;
    assign layer_1_weights[24][109] = 6'sd3;
    assign layer_1_weights[24][110] = -6'sd2;
    assign layer_1_weights[24][111] = 6'sd2;
    assign layer_1_weights[24][112] = 6'sd5;
    assign layer_1_weights[24][113] = 6'sd3;
    assign layer_1_weights[24][114] = 6'sd0;
    assign layer_1_weights[24][115] = 6'sd0;
    assign layer_1_weights[24][116] = 6'sd1;
    assign layer_1_weights[24][117] = 6'sd1;
    assign layer_1_weights[24][118] = 6'sd0;
    assign layer_1_weights[24][119] = 6'sd2;
    assign layer_1_weights[24][120] = -6'sd2;
    assign layer_1_weights[24][121] = 6'sd3;
    assign layer_1_weights[24][122] = -6'sd4;
    assign layer_1_weights[24][123] = 6'sd0;
    assign layer_1_weights[24][124] = 6'sd4;
    assign layer_1_weights[24][125] = -6'sd2;
    assign layer_1_weights[24][126] = 6'sd0;
    assign layer_1_weights[24][127] = 6'sd0;
    assign layer_1_weights[24][128] = 6'sd0;
    assign layer_1_weights[24][129] = 6'sd2;
    assign layer_1_weights[24][130] = 6'sd4;
    assign layer_1_weights[24][131] = -6'sd6;
    assign layer_1_weights[24][132] = 6'sd1;
    assign layer_1_weights[24][133] = 6'sd1;
    assign layer_1_weights[24][134] = -6'sd12;
    assign layer_1_weights[24][135] = -6'sd5;
    assign layer_1_weights[24][136] = 6'sd1;
    assign layer_1_weights[24][137] = 6'sd1;
    assign layer_1_weights[24][138] = -6'sd1;
    assign layer_1_weights[24][139] = -6'sd5;
    assign layer_1_weights[24][140] = -6'sd7;
    assign layer_1_weights[24][141] = -6'sd9;
    assign layer_1_weights[24][142] = -6'sd1;
    assign layer_1_weights[24][143] = -6'sd1;
    assign layer_1_biases[24] = -6'sd3;
    assign layer_1_weights[25][0] = 6'sd2;
    assign layer_1_weights[25][1] = -6'sd1;
    assign layer_1_weights[25][2] = 6'sd1;
    assign layer_1_weights[25][3] = -6'sd2;
    assign layer_1_weights[25][4] = 6'sd7;
    assign layer_1_weights[25][5] = -6'sd2;
    assign layer_1_weights[25][6] = -6'sd4;
    assign layer_1_weights[25][7] = 6'sd3;
    assign layer_1_weights[25][8] = 6'sd7;
    assign layer_1_weights[25][9] = 6'sd6;
    assign layer_1_weights[25][10] = 6'sd0;
    assign layer_1_weights[25][11] = 6'sd1;
    assign layer_1_weights[25][12] = 6'sd0;
    assign layer_1_weights[25][13] = 6'sd0;
    assign layer_1_weights[25][14] = 6'sd4;
    assign layer_1_weights[25][15] = -6'sd3;
    assign layer_1_weights[25][16] = -6'sd5;
    assign layer_1_weights[25][17] = -6'sd8;
    assign layer_1_weights[25][18] = -6'sd7;
    assign layer_1_weights[25][19] = -6'sd1;
    assign layer_1_weights[25][20] = -6'sd11;
    assign layer_1_weights[25][21] = -6'sd8;
    assign layer_1_weights[25][22] = -6'sd5;
    assign layer_1_weights[25][23] = 6'sd0;
    assign layer_1_weights[25][24] = 6'sd1;
    assign layer_1_weights[25][25] = 6'sd6;
    assign layer_1_weights[25][26] = 6'sd2;
    assign layer_1_weights[25][27] = -6'sd3;
    assign layer_1_weights[25][28] = -6'sd3;
    assign layer_1_weights[25][29] = -6'sd1;
    assign layer_1_weights[25][30] = -6'sd5;
    assign layer_1_weights[25][31] = -6'sd5;
    assign layer_1_weights[25][32] = -6'sd4;
    assign layer_1_weights[25][33] = -6'sd4;
    assign layer_1_weights[25][34] = -6'sd4;
    assign layer_1_weights[25][35] = -6'sd5;
    assign layer_1_weights[25][36] = -6'sd2;
    assign layer_1_weights[25][37] = 6'sd3;
    assign layer_1_weights[25][38] = -6'sd1;
    assign layer_1_weights[25][39] = -6'sd2;
    assign layer_1_weights[25][40] = -6'sd5;
    assign layer_1_weights[25][41] = -6'sd7;
    assign layer_1_weights[25][42] = 6'sd1;
    assign layer_1_weights[25][43] = 6'sd6;
    assign layer_1_weights[25][44] = 6'sd8;
    assign layer_1_weights[25][45] = 6'sd7;
    assign layer_1_weights[25][46] = 6'sd6;
    assign layer_1_weights[25][47] = 6'sd0;
    assign layer_1_weights[25][48] = 6'sd7;
    assign layer_1_weights[25][49] = 6'sd4;
    assign layer_1_weights[25][50] = -6'sd2;
    assign layer_1_weights[25][51] = 6'sd0;
    assign layer_1_weights[25][52] = -6'sd3;
    assign layer_1_weights[25][53] = 6'sd0;
    assign layer_1_weights[25][54] = 6'sd5;
    assign layer_1_weights[25][55] = 6'sd6;
    assign layer_1_weights[25][56] = 6'sd9;
    assign layer_1_weights[25][57] = 6'sd8;
    assign layer_1_weights[25][58] = 6'sd7;
    assign layer_1_weights[25][59] = 6'sd3;
    assign layer_1_weights[25][60] = 6'sd3;
    assign layer_1_weights[25][61] = -6'sd2;
    assign layer_1_weights[25][62] = -6'sd2;
    assign layer_1_weights[25][63] = 6'sd2;
    assign layer_1_weights[25][64] = 6'sd2;
    assign layer_1_weights[25][65] = 6'sd1;
    assign layer_1_weights[25][66] = -6'sd4;
    assign layer_1_weights[25][67] = -6'sd9;
    assign layer_1_weights[25][68] = -6'sd10;
    assign layer_1_weights[25][69] = -6'sd4;
    assign layer_1_weights[25][70] = -6'sd2;
    assign layer_1_weights[25][71] = 6'sd7;
    assign layer_1_weights[25][72] = 6'sd1;
    assign layer_1_weights[25][73] = -6'sd1;
    assign layer_1_weights[25][74] = -6'sd1;
    assign layer_1_weights[25][75] = 6'sd0;
    assign layer_1_weights[25][76] = 6'sd1;
    assign layer_1_weights[25][77] = 6'sd5;
    assign layer_1_weights[25][78] = -6'sd2;
    assign layer_1_weights[25][79] = -6'sd1;
    assign layer_1_weights[25][80] = -6'sd4;
    assign layer_1_weights[25][81] = -6'sd3;
    assign layer_1_weights[25][82] = -6'sd4;
    assign layer_1_weights[25][83] = -6'sd3;
    assign layer_1_weights[25][84] = 6'sd1;
    assign layer_1_weights[25][85] = -6'sd4;
    assign layer_1_weights[25][86] = 6'sd2;
    assign layer_1_weights[25][87] = 6'sd2;
    assign layer_1_weights[25][88] = 6'sd3;
    assign layer_1_weights[25][89] = 6'sd1;
    assign layer_1_weights[25][90] = -6'sd1;
    assign layer_1_weights[25][91] = 6'sd0;
    assign layer_1_weights[25][92] = 6'sd0;
    assign layer_1_weights[25][93] = -6'sd3;
    assign layer_1_weights[25][94] = -6'sd2;
    assign layer_1_weights[25][95] = 6'sd4;
    assign layer_1_weights[25][96] = 6'sd0;
    assign layer_1_weights[25][97] = -6'sd6;
    assign layer_1_weights[25][98] = 6'sd1;
    assign layer_1_weights[25][99] = 6'sd2;
    assign layer_1_weights[25][100] = 6'sd3;
    assign layer_1_weights[25][101] = 6'sd4;
    assign layer_1_weights[25][102] = -6'sd2;
    assign layer_1_weights[25][103] = -6'sd3;
    assign layer_1_weights[25][104] = 6'sd0;
    assign layer_1_weights[25][105] = -6'sd3;
    assign layer_1_weights[25][106] = -6'sd5;
    assign layer_1_weights[25][107] = 6'sd6;
    assign layer_1_weights[25][108] = -6'sd1;
    assign layer_1_weights[25][109] = -6'sd8;
    assign layer_1_weights[25][110] = 6'sd0;
    assign layer_1_weights[25][111] = 6'sd0;
    assign layer_1_weights[25][112] = -6'sd2;
    assign layer_1_weights[25][113] = -6'sd1;
    assign layer_1_weights[25][114] = -6'sd4;
    assign layer_1_weights[25][115] = -6'sd2;
    assign layer_1_weights[25][116] = -6'sd1;
    assign layer_1_weights[25][117] = -6'sd2;
    assign layer_1_weights[25][118] = 6'sd3;
    assign layer_1_weights[25][119] = -6'sd5;
    assign layer_1_weights[25][120] = 6'sd0;
    assign layer_1_weights[25][121] = -6'sd8;
    assign layer_1_weights[25][122] = -6'sd2;
    assign layer_1_weights[25][123] = 6'sd0;
    assign layer_1_weights[25][124] = 6'sd5;
    assign layer_1_weights[25][125] = 6'sd0;
    assign layer_1_weights[25][126] = 6'sd1;
    assign layer_1_weights[25][127] = -6'sd2;
    assign layer_1_weights[25][128] = 6'sd1;
    assign layer_1_weights[25][129] = -6'sd5;
    assign layer_1_weights[25][130] = -6'sd5;
    assign layer_1_weights[25][131] = 6'sd1;
    assign layer_1_weights[25][132] = -6'sd1;
    assign layer_1_weights[25][133] = 6'sd5;
    assign layer_1_weights[25][134] = -6'sd2;
    assign layer_1_weights[25][135] = -6'sd10;
    assign layer_1_weights[25][136] = 6'sd0;
    assign layer_1_weights[25][137] = 6'sd1;
    assign layer_1_weights[25][138] = -6'sd6;
    assign layer_1_weights[25][139] = 6'sd6;
    assign layer_1_weights[25][140] = 6'sd0;
    assign layer_1_weights[25][141] = 6'sd4;
    assign layer_1_weights[25][142] = -6'sd2;
    assign layer_1_weights[25][143] = -6'sd2;
    assign layer_1_biases[25] = 6'sd6;
    assign layer_1_weights[26][0] = 6'sd2;
    assign layer_1_weights[26][1] = 6'sd1;
    assign layer_1_weights[26][2] = -6'sd3;
    assign layer_1_weights[26][3] = -6'sd4;
    assign layer_1_weights[26][4] = -6'sd7;
    assign layer_1_weights[26][5] = -6'sd7;
    assign layer_1_weights[26][6] = -6'sd2;
    assign layer_1_weights[26][7] = -6'sd4;
    assign layer_1_weights[26][8] = -6'sd14;
    assign layer_1_weights[26][9] = -6'sd11;
    assign layer_1_weights[26][10] = 6'sd2;
    assign layer_1_weights[26][11] = -6'sd2;
    assign layer_1_weights[26][12] = 6'sd0;
    assign layer_1_weights[26][13] = -6'sd1;
    assign layer_1_weights[26][14] = -6'sd2;
    assign layer_1_weights[26][15] = -6'sd10;
    assign layer_1_weights[26][16] = -6'sd7;
    assign layer_1_weights[26][17] = -6'sd6;
    assign layer_1_weights[26][18] = -6'sd6;
    assign layer_1_weights[26][19] = -6'sd4;
    assign layer_1_weights[26][20] = -6'sd4;
    assign layer_1_weights[26][21] = -6'sd7;
    assign layer_1_weights[26][22] = 6'sd0;
    assign layer_1_weights[26][23] = -6'sd1;
    assign layer_1_weights[26][24] = 6'sd0;
    assign layer_1_weights[26][25] = 6'sd2;
    assign layer_1_weights[26][26] = -6'sd7;
    assign layer_1_weights[26][27] = -6'sd5;
    assign layer_1_weights[26][28] = -6'sd1;
    assign layer_1_weights[26][29] = 6'sd2;
    assign layer_1_weights[26][30] = -6'sd1;
    assign layer_1_weights[26][31] = 6'sd1;
    assign layer_1_weights[26][32] = 6'sd2;
    assign layer_1_weights[26][33] = -6'sd1;
    assign layer_1_weights[26][34] = -6'sd1;
    assign layer_1_weights[26][35] = 6'sd2;
    assign layer_1_weights[26][36] = 6'sd8;
    assign layer_1_weights[26][37] = 6'sd0;
    assign layer_1_weights[26][38] = 6'sd2;
    assign layer_1_weights[26][39] = -6'sd2;
    assign layer_1_weights[26][40] = 6'sd1;
    assign layer_1_weights[26][41] = 6'sd1;
    assign layer_1_weights[26][42] = 6'sd3;
    assign layer_1_weights[26][43] = 6'sd5;
    assign layer_1_weights[26][44] = 6'sd4;
    assign layer_1_weights[26][45] = 6'sd3;
    assign layer_1_weights[26][46] = 6'sd5;
    assign layer_1_weights[26][47] = 6'sd2;
    assign layer_1_weights[26][48] = 6'sd5;
    assign layer_1_weights[26][49] = -6'sd2;
    assign layer_1_weights[26][50] = 6'sd1;
    assign layer_1_weights[26][51] = 6'sd1;
    assign layer_1_weights[26][52] = 6'sd4;
    assign layer_1_weights[26][53] = 6'sd7;
    assign layer_1_weights[26][54] = 6'sd5;
    assign layer_1_weights[26][55] = 6'sd3;
    assign layer_1_weights[26][56] = 6'sd3;
    assign layer_1_weights[26][57] = 6'sd5;
    assign layer_1_weights[26][58] = 6'sd5;
    assign layer_1_weights[26][59] = 6'sd0;
    assign layer_1_weights[26][60] = 6'sd12;
    assign layer_1_weights[26][61] = 6'sd0;
    assign layer_1_weights[26][62] = -6'sd2;
    assign layer_1_weights[26][63] = 6'sd3;
    assign layer_1_weights[26][64] = 6'sd2;
    assign layer_1_weights[26][65] = 6'sd2;
    assign layer_1_weights[26][66] = 6'sd3;
    assign layer_1_weights[26][67] = 6'sd2;
    assign layer_1_weights[26][68] = 6'sd2;
    assign layer_1_weights[26][69] = -6'sd3;
    assign layer_1_weights[26][70] = -6'sd4;
    assign layer_1_weights[26][71] = 6'sd6;
    assign layer_1_weights[26][72] = 6'sd6;
    assign layer_1_weights[26][73] = 6'sd1;
    assign layer_1_weights[26][74] = 6'sd0;
    assign layer_1_weights[26][75] = -6'sd3;
    assign layer_1_weights[26][76] = -6'sd6;
    assign layer_1_weights[26][77] = -6'sd3;
    assign layer_1_weights[26][78] = 6'sd2;
    assign layer_1_weights[26][79] = 6'sd3;
    assign layer_1_weights[26][80] = 6'sd3;
    assign layer_1_weights[26][81] = -6'sd3;
    assign layer_1_weights[26][82] = 6'sd1;
    assign layer_1_weights[26][83] = 6'sd4;
    assign layer_1_weights[26][84] = 6'sd8;
    assign layer_1_weights[26][85] = 6'sd1;
    assign layer_1_weights[26][86] = 6'sd2;
    assign layer_1_weights[26][87] = 6'sd1;
    assign layer_1_weights[26][88] = -6'sd2;
    assign layer_1_weights[26][89] = -6'sd3;
    assign layer_1_weights[26][90] = 6'sd0;
    assign layer_1_weights[26][91] = 6'sd3;
    assign layer_1_weights[26][92] = 6'sd0;
    assign layer_1_weights[26][93] = 6'sd4;
    assign layer_1_weights[26][94] = 6'sd0;
    assign layer_1_weights[26][95] = -6'sd2;
    assign layer_1_weights[26][96] = -6'sd6;
    assign layer_1_weights[26][97] = 6'sd2;
    assign layer_1_weights[26][98] = 6'sd0;
    assign layer_1_weights[26][99] = -6'sd2;
    assign layer_1_weights[26][100] = -6'sd4;
    assign layer_1_weights[26][101] = -6'sd5;
    assign layer_1_weights[26][102] = -6'sd3;
    assign layer_1_weights[26][103] = 6'sd1;
    assign layer_1_weights[26][104] = 6'sd0;
    assign layer_1_weights[26][105] = 6'sd2;
    assign layer_1_weights[26][106] = 6'sd0;
    assign layer_1_weights[26][107] = 6'sd1;
    assign layer_1_weights[26][108] = 6'sd4;
    assign layer_1_weights[26][109] = 6'sd2;
    assign layer_1_weights[26][110] = 6'sd2;
    assign layer_1_weights[26][111] = -6'sd1;
    assign layer_1_weights[26][112] = -6'sd3;
    assign layer_1_weights[26][113] = -6'sd2;
    assign layer_1_weights[26][114] = 6'sd1;
    assign layer_1_weights[26][115] = 6'sd2;
    assign layer_1_weights[26][116] = -6'sd2;
    assign layer_1_weights[26][117] = -6'sd7;
    assign layer_1_weights[26][118] = -6'sd6;
    assign layer_1_weights[26][119] = -6'sd2;
    assign layer_1_weights[26][120] = 6'sd2;
    assign layer_1_weights[26][121] = 6'sd8;
    assign layer_1_weights[26][122] = 6'sd4;
    assign layer_1_weights[26][123] = 6'sd1;
    assign layer_1_weights[26][124] = 6'sd1;
    assign layer_1_weights[26][125] = -6'sd1;
    assign layer_1_weights[26][126] = 6'sd1;
    assign layer_1_weights[26][127] = -6'sd1;
    assign layer_1_weights[26][128] = 6'sd0;
    assign layer_1_weights[26][129] = 6'sd1;
    assign layer_1_weights[26][130] = -6'sd3;
    assign layer_1_weights[26][131] = -6'sd6;
    assign layer_1_weights[26][132] = 6'sd0;
    assign layer_1_weights[26][133] = 6'sd1;
    assign layer_1_weights[26][134] = 6'sd5;
    assign layer_1_weights[26][135] = 6'sd10;
    assign layer_1_weights[26][136] = 6'sd11;
    assign layer_1_weights[26][137] = 6'sd8;
    assign layer_1_weights[26][138] = 6'sd7;
    assign layer_1_weights[26][139] = 6'sd6;
    assign layer_1_weights[26][140] = 6'sd7;
    assign layer_1_weights[26][141] = 6'sd1;
    assign layer_1_weights[26][142] = -6'sd1;
    assign layer_1_weights[26][143] = 6'sd1;
    assign layer_1_biases[26] = 6'sd2;
    assign layer_1_weights[27][0] = -6'sd1;
    assign layer_1_weights[27][1] = 6'sd0;
    assign layer_1_weights[27][2] = 6'sd1;
    assign layer_1_weights[27][3] = 6'sd0;
    assign layer_1_weights[27][4] = 6'sd6;
    assign layer_1_weights[27][5] = -6'sd8;
    assign layer_1_weights[27][6] = 6'sd2;
    assign layer_1_weights[27][7] = 6'sd7;
    assign layer_1_weights[27][8] = -6'sd3;
    assign layer_1_weights[27][9] = -6'sd2;
    assign layer_1_weights[27][10] = -6'sd1;
    assign layer_1_weights[27][11] = 6'sd2;
    assign layer_1_weights[27][12] = 6'sd0;
    assign layer_1_weights[27][13] = -6'sd1;
    assign layer_1_weights[27][14] = 6'sd0;
    assign layer_1_weights[27][15] = 6'sd1;
    assign layer_1_weights[27][16] = 6'sd4;
    assign layer_1_weights[27][17] = 6'sd3;
    assign layer_1_weights[27][18] = -6'sd6;
    assign layer_1_weights[27][19] = 6'sd0;
    assign layer_1_weights[27][20] = -6'sd3;
    assign layer_1_weights[27][21] = -6'sd4;
    assign layer_1_weights[27][22] = 6'sd6;
    assign layer_1_weights[27][23] = 6'sd2;
    assign layer_1_weights[27][24] = 6'sd0;
    assign layer_1_weights[27][25] = 6'sd5;
    assign layer_1_weights[27][26] = 6'sd6;
    assign layer_1_weights[27][27] = 6'sd7;
    assign layer_1_weights[27][28] = 6'sd3;
    assign layer_1_weights[27][29] = 6'sd3;
    assign layer_1_weights[27][30] = -6'sd3;
    assign layer_1_weights[27][31] = -6'sd3;
    assign layer_1_weights[27][32] = -6'sd2;
    assign layer_1_weights[27][33] = -6'sd2;
    assign layer_1_weights[27][34] = 6'sd3;
    assign layer_1_weights[27][35] = 6'sd8;
    assign layer_1_weights[27][36] = 6'sd4;
    assign layer_1_weights[27][37] = 6'sd6;
    assign layer_1_weights[27][38] = -6'sd3;
    assign layer_1_weights[27][39] = 6'sd1;
    assign layer_1_weights[27][40] = 6'sd6;
    assign layer_1_weights[27][41] = 6'sd2;
    assign layer_1_weights[27][42] = -6'sd5;
    assign layer_1_weights[27][43] = 6'sd0;
    assign layer_1_weights[27][44] = 6'sd2;
    assign layer_1_weights[27][45] = 6'sd4;
    assign layer_1_weights[27][46] = 6'sd7;
    assign layer_1_weights[27][47] = 6'sd5;
    assign layer_1_weights[27][48] = -6'sd2;
    assign layer_1_weights[27][49] = 6'sd4;
    assign layer_1_weights[27][50] = -6'sd1;
    assign layer_1_weights[27][51] = -6'sd1;
    assign layer_1_weights[27][52] = 6'sd2;
    assign layer_1_weights[27][53] = 6'sd4;
    assign layer_1_weights[27][54] = -6'sd2;
    assign layer_1_weights[27][55] = 6'sd6;
    assign layer_1_weights[27][56] = 6'sd3;
    assign layer_1_weights[27][57] = 6'sd4;
    assign layer_1_weights[27][58] = 6'sd4;
    assign layer_1_weights[27][59] = 6'sd0;
    assign layer_1_weights[27][60] = 6'sd11;
    assign layer_1_weights[27][61] = -6'sd10;
    assign layer_1_weights[27][62] = -6'sd5;
    assign layer_1_weights[27][63] = -6'sd1;
    assign layer_1_weights[27][64] = 6'sd3;
    assign layer_1_weights[27][65] = -6'sd1;
    assign layer_1_weights[27][66] = -6'sd2;
    assign layer_1_weights[27][67] = 6'sd4;
    assign layer_1_weights[27][68] = -6'sd2;
    assign layer_1_weights[27][69] = -6'sd2;
    assign layer_1_weights[27][70] = -6'sd1;
    assign layer_1_weights[27][71] = 6'sd3;
    assign layer_1_weights[27][72] = 6'sd6;
    assign layer_1_weights[27][73] = -6'sd2;
    assign layer_1_weights[27][74] = -6'sd4;
    assign layer_1_weights[27][75] = 6'sd2;
    assign layer_1_weights[27][76] = -6'sd1;
    assign layer_1_weights[27][77] = -6'sd4;
    assign layer_1_weights[27][78] = 6'sd1;
    assign layer_1_weights[27][79] = -6'sd3;
    assign layer_1_weights[27][80] = 6'sd2;
    assign layer_1_weights[27][81] = 6'sd1;
    assign layer_1_weights[27][82] = 6'sd0;
    assign layer_1_weights[27][83] = -6'sd3;
    assign layer_1_weights[27][84] = 6'sd3;
    assign layer_1_weights[27][85] = 6'sd6;
    assign layer_1_weights[27][86] = 6'sd4;
    assign layer_1_weights[27][87] = 6'sd2;
    assign layer_1_weights[27][88] = 6'sd0;
    assign layer_1_weights[27][89] = 6'sd0;
    assign layer_1_weights[27][90] = 6'sd0;
    assign layer_1_weights[27][91] = -6'sd5;
    assign layer_1_weights[27][92] = 6'sd1;
    assign layer_1_weights[27][93] = 6'sd2;
    assign layer_1_weights[27][94] = -6'sd1;
    assign layer_1_weights[27][95] = 6'sd4;
    assign layer_1_weights[27][96] = 6'sd0;
    assign layer_1_weights[27][97] = 6'sd8;
    assign layer_1_weights[27][98] = 6'sd0;
    assign layer_1_weights[27][99] = -6'sd1;
    assign layer_1_weights[27][100] = 6'sd3;
    assign layer_1_weights[27][101] = 6'sd3;
    assign layer_1_weights[27][102] = -6'sd2;
    assign layer_1_weights[27][103] = -6'sd5;
    assign layer_1_weights[27][104] = -6'sd2;
    assign layer_1_weights[27][105] = 6'sd0;
    assign layer_1_weights[27][106] = -6'sd4;
    assign layer_1_weights[27][107] = -6'sd1;
    assign layer_1_weights[27][108] = -6'sd1;
    assign layer_1_weights[27][109] = -6'sd6;
    assign layer_1_weights[27][110] = -6'sd5;
    assign layer_1_weights[27][111] = -6'sd2;
    assign layer_1_weights[27][112] = 6'sd3;
    assign layer_1_weights[27][113] = 6'sd2;
    assign layer_1_weights[27][114] = 6'sd0;
    assign layer_1_weights[27][115] = -6'sd1;
    assign layer_1_weights[27][116] = -6'sd3;
    assign layer_1_weights[27][117] = -6'sd2;
    assign layer_1_weights[27][118] = -6'sd2;
    assign layer_1_weights[27][119] = -6'sd3;
    assign layer_1_weights[27][120] = -6'sd1;
    assign layer_1_weights[27][121] = 6'sd4;
    assign layer_1_weights[27][122] = 6'sd0;
    assign layer_1_weights[27][123] = -6'sd2;
    assign layer_1_weights[27][124] = 6'sd0;
    assign layer_1_weights[27][125] = 6'sd5;
    assign layer_1_weights[27][126] = 6'sd2;
    assign layer_1_weights[27][127] = 6'sd0;
    assign layer_1_weights[27][128] = -6'sd2;
    assign layer_1_weights[27][129] = -6'sd7;
    assign layer_1_weights[27][130] = -6'sd12;
    assign layer_1_weights[27][131] = -6'sd2;
    assign layer_1_weights[27][132] = 6'sd0;
    assign layer_1_weights[27][133] = -6'sd2;
    assign layer_1_weights[27][134] = 6'sd0;
    assign layer_1_weights[27][135] = 6'sd1;
    assign layer_1_weights[27][136] = 6'sd0;
    assign layer_1_weights[27][137] = 6'sd4;
    assign layer_1_weights[27][138] = 6'sd0;
    assign layer_1_weights[27][139] = 6'sd4;
    assign layer_1_weights[27][140] = 6'sd7;
    assign layer_1_weights[27][141] = -6'sd2;
    assign layer_1_weights[27][142] = 6'sd0;
    assign layer_1_weights[27][143] = 6'sd1;
    assign layer_1_biases[27] = 6'sd1;
    assign layer_1_weights[28][0] = 6'sd0;
    assign layer_1_weights[28][1] = -6'sd1;
    assign layer_1_weights[28][2] = -6'sd1;
    assign layer_1_weights[28][3] = -6'sd1;
    assign layer_1_weights[28][4] = 6'sd2;
    assign layer_1_weights[28][5] = 6'sd5;
    assign layer_1_weights[28][6] = 6'sd4;
    assign layer_1_weights[28][7] = 6'sd0;
    assign layer_1_weights[28][8] = 6'sd2;
    assign layer_1_weights[28][9] = -6'sd5;
    assign layer_1_weights[28][10] = 6'sd0;
    assign layer_1_weights[28][11] = -6'sd1;
    assign layer_1_weights[28][12] = 6'sd1;
    assign layer_1_weights[28][13] = -6'sd1;
    assign layer_1_weights[28][14] = 6'sd3;
    assign layer_1_weights[28][15] = 6'sd3;
    assign layer_1_weights[28][16] = 6'sd4;
    assign layer_1_weights[28][17] = 6'sd1;
    assign layer_1_weights[28][18] = -6'sd1;
    assign layer_1_weights[28][19] = 6'sd2;
    assign layer_1_weights[28][20] = 6'sd2;
    assign layer_1_weights[28][21] = -6'sd1;
    assign layer_1_weights[28][22] = -6'sd4;
    assign layer_1_weights[28][23] = 6'sd1;
    assign layer_1_weights[28][24] = 6'sd1;
    assign layer_1_weights[28][25] = -6'sd2;
    assign layer_1_weights[28][26] = -6'sd6;
    assign layer_1_weights[28][27] = -6'sd2;
    assign layer_1_weights[28][28] = -6'sd6;
    assign layer_1_weights[28][29] = 6'sd0;
    assign layer_1_weights[28][30] = 6'sd2;
    assign layer_1_weights[28][31] = 6'sd1;
    assign layer_1_weights[28][32] = 6'sd1;
    assign layer_1_weights[28][33] = 6'sd2;
    assign layer_1_weights[28][34] = 6'sd2;
    assign layer_1_weights[28][35] = 6'sd1;
    assign layer_1_weights[28][36] = 6'sd5;
    assign layer_1_weights[28][37] = 6'sd9;
    assign layer_1_weights[28][38] = 6'sd0;
    assign layer_1_weights[28][39] = 6'sd2;
    assign layer_1_weights[28][40] = -6'sd6;
    assign layer_1_weights[28][41] = -6'sd5;
    assign layer_1_weights[28][42] = 6'sd1;
    assign layer_1_weights[28][43] = 6'sd1;
    assign layer_1_weights[28][44] = 6'sd1;
    assign layer_1_weights[28][45] = 6'sd2;
    assign layer_1_weights[28][46] = 6'sd2;
    assign layer_1_weights[28][47] = 6'sd2;
    assign layer_1_weights[28][48] = 6'sd1;
    assign layer_1_weights[28][49] = 6'sd10;
    assign layer_1_weights[28][50] = 6'sd8;
    assign layer_1_weights[28][51] = 6'sd7;
    assign layer_1_weights[28][52] = -6'sd1;
    assign layer_1_weights[28][53] = -6'sd2;
    assign layer_1_weights[28][54] = 6'sd2;
    assign layer_1_weights[28][55] = 6'sd4;
    assign layer_1_weights[28][56] = 6'sd4;
    assign layer_1_weights[28][57] = 6'sd2;
    assign layer_1_weights[28][58] = -6'sd2;
    assign layer_1_weights[28][59] = -6'sd1;
    assign layer_1_weights[28][60] = 6'sd1;
    assign layer_1_weights[28][61] = 6'sd2;
    assign layer_1_weights[28][62] = 6'sd2;
    assign layer_1_weights[28][63] = 6'sd1;
    assign layer_1_weights[28][64] = -6'sd5;
    assign layer_1_weights[28][65] = 6'sd1;
    assign layer_1_weights[28][66] = 6'sd1;
    assign layer_1_weights[28][67] = -6'sd1;
    assign layer_1_weights[28][68] = 6'sd1;
    assign layer_1_weights[28][69] = -6'sd2;
    assign layer_1_weights[28][70] = -6'sd2;
    assign layer_1_weights[28][71] = 6'sd4;
    assign layer_1_weights[28][72] = 6'sd5;
    assign layer_1_weights[28][73] = -6'sd7;
    assign layer_1_weights[28][74] = -6'sd8;
    assign layer_1_weights[28][75] = -6'sd7;
    assign layer_1_weights[28][76] = -6'sd4;
    assign layer_1_weights[28][77] = 6'sd7;
    assign layer_1_weights[28][78] = 6'sd5;
    assign layer_1_weights[28][79] = 6'sd0;
    assign layer_1_weights[28][80] = -6'sd5;
    assign layer_1_weights[28][81] = -6'sd7;
    assign layer_1_weights[28][82] = -6'sd1;
    assign layer_1_weights[28][83] = -6'sd1;
    assign layer_1_weights[28][84] = 6'sd4;
    assign layer_1_weights[28][85] = -6'sd4;
    assign layer_1_weights[28][86] = -6'sd8;
    assign layer_1_weights[28][87] = -6'sd5;
    assign layer_1_weights[28][88] = 6'sd3;
    assign layer_1_weights[28][89] = 6'sd7;
    assign layer_1_weights[28][90] = 6'sd2;
    assign layer_1_weights[28][91] = -6'sd2;
    assign layer_1_weights[28][92] = 6'sd0;
    assign layer_1_weights[28][93] = 6'sd0;
    assign layer_1_weights[28][94] = 6'sd2;
    assign layer_1_weights[28][95] = 6'sd3;
    assign layer_1_weights[28][96] = -6'sd1;
    assign layer_1_weights[28][97] = 6'sd2;
    assign layer_1_weights[28][98] = 6'sd0;
    assign layer_1_weights[28][99] = 6'sd5;
    assign layer_1_weights[28][100] = 6'sd5;
    assign layer_1_weights[28][101] = 6'sd1;
    assign layer_1_weights[28][102] = -6'sd3;
    assign layer_1_weights[28][103] = 6'sd1;
    assign layer_1_weights[28][104] = 6'sd2;
    assign layer_1_weights[28][105] = 6'sd0;
    assign layer_1_weights[28][106] = 6'sd4;
    assign layer_1_weights[28][107] = 6'sd5;
    assign layer_1_weights[28][108] = 6'sd11;
    assign layer_1_weights[28][109] = 6'sd4;
    assign layer_1_weights[28][110] = 6'sd4;
    assign layer_1_weights[28][111] = 6'sd4;
    assign layer_1_weights[28][112] = 6'sd1;
    assign layer_1_weights[28][113] = -6'sd1;
    assign layer_1_weights[28][114] = -6'sd1;
    assign layer_1_weights[28][115] = 6'sd0;
    assign layer_1_weights[28][116] = 6'sd2;
    assign layer_1_weights[28][117] = 6'sd1;
    assign layer_1_weights[28][118] = 6'sd4;
    assign layer_1_weights[28][119] = -6'sd4;
    assign layer_1_weights[28][120] = 6'sd1;
    assign layer_1_weights[28][121] = -6'sd5;
    assign layer_1_weights[28][122] = 6'sd2;
    assign layer_1_weights[28][123] = 6'sd1;
    assign layer_1_weights[28][124] = 6'sd2;
    assign layer_1_weights[28][125] = 6'sd2;
    assign layer_1_weights[28][126] = 6'sd1;
    assign layer_1_weights[28][127] = -6'sd1;
    assign layer_1_weights[28][128] = 6'sd0;
    assign layer_1_weights[28][129] = -6'sd1;
    assign layer_1_weights[28][130] = -6'sd2;
    assign layer_1_weights[28][131] = 6'sd6;
    assign layer_1_weights[28][132] = 6'sd0;
    assign layer_1_weights[28][133] = -6'sd4;
    assign layer_1_weights[28][134] = -6'sd2;
    assign layer_1_weights[28][135] = -6'sd2;
    assign layer_1_weights[28][136] = 6'sd1;
    assign layer_1_weights[28][137] = -6'sd6;
    assign layer_1_weights[28][138] = 6'sd1;
    assign layer_1_weights[28][139] = -6'sd4;
    assign layer_1_weights[28][140] = -6'sd2;
    assign layer_1_weights[28][141] = -6'sd10;
    assign layer_1_weights[28][142] = 6'sd1;
    assign layer_1_weights[28][143] = 6'sd2;
    assign layer_1_biases[28] = -6'sd1;
    assign layer_1_weights[29][0] = -6'sd2;
    assign layer_1_weights[29][1] = -6'sd2;
    assign layer_1_weights[29][2] = 6'sd5;
    assign layer_1_weights[29][3] = 6'sd8;
    assign layer_1_weights[29][4] = 6'sd8;
    assign layer_1_weights[29][5] = 6'sd2;
    assign layer_1_weights[29][6] = -6'sd4;
    assign layer_1_weights[29][7] = 6'sd10;
    assign layer_1_weights[29][8] = 6'sd8;
    assign layer_1_weights[29][9] = 6'sd11;
    assign layer_1_weights[29][10] = -6'sd2;
    assign layer_1_weights[29][11] = 6'sd0;
    assign layer_1_weights[29][12] = -6'sd2;
    assign layer_1_weights[29][13] = 6'sd1;
    assign layer_1_weights[29][14] = 6'sd6;
    assign layer_1_weights[29][15] = 6'sd7;
    assign layer_1_weights[29][16] = 6'sd8;
    assign layer_1_weights[29][17] = 6'sd0;
    assign layer_1_weights[29][18] = 6'sd2;
    assign layer_1_weights[29][19] = -6'sd2;
    assign layer_1_weights[29][20] = 6'sd5;
    assign layer_1_weights[29][21] = -6'sd2;
    assign layer_1_weights[29][22] = 6'sd2;
    assign layer_1_weights[29][23] = 6'sd2;
    assign layer_1_weights[29][24] = 6'sd0;
    assign layer_1_weights[29][25] = 6'sd0;
    assign layer_1_weights[29][26] = 6'sd4;
    assign layer_1_weights[29][27] = -6'sd2;
    assign layer_1_weights[29][28] = -6'sd4;
    assign layer_1_weights[29][29] = 6'sd1;
    assign layer_1_weights[29][30] = 6'sd2;
    assign layer_1_weights[29][31] = -6'sd1;
    assign layer_1_weights[29][32] = 6'sd0;
    assign layer_1_weights[29][33] = -6'sd2;
    assign layer_1_weights[29][34] = -6'sd1;
    assign layer_1_weights[29][35] = 6'sd7;
    assign layer_1_weights[29][36] = -6'sd1;
    assign layer_1_weights[29][37] = 6'sd8;
    assign layer_1_weights[29][38] = -6'sd3;
    assign layer_1_weights[29][39] = 6'sd0;
    assign layer_1_weights[29][40] = -6'sd4;
    assign layer_1_weights[29][41] = 6'sd1;
    assign layer_1_weights[29][42] = -6'sd5;
    assign layer_1_weights[29][43] = -6'sd7;
    assign layer_1_weights[29][44] = -6'sd2;
    assign layer_1_weights[29][45] = 6'sd0;
    assign layer_1_weights[29][46] = -6'sd7;
    assign layer_1_weights[29][47] = -6'sd1;
    assign layer_1_weights[29][48] = -6'sd2;
    assign layer_1_weights[29][49] = 6'sd5;
    assign layer_1_weights[29][50] = -6'sd2;
    assign layer_1_weights[29][51] = -6'sd4;
    assign layer_1_weights[29][52] = -6'sd1;
    assign layer_1_weights[29][53] = 6'sd1;
    assign layer_1_weights[29][54] = 6'sd1;
    assign layer_1_weights[29][55] = 6'sd1;
    assign layer_1_weights[29][56] = -6'sd3;
    assign layer_1_weights[29][57] = -6'sd3;
    assign layer_1_weights[29][58] = -6'sd4;
    assign layer_1_weights[29][59] = -6'sd5;
    assign layer_1_weights[29][60] = -6'sd4;
    assign layer_1_weights[29][61] = -6'sd8;
    assign layer_1_weights[29][62] = 6'sd1;
    assign layer_1_weights[29][63] = 6'sd0;
    assign layer_1_weights[29][64] = 6'sd1;
    assign layer_1_weights[29][65] = 6'sd2;
    assign layer_1_weights[29][66] = 6'sd5;
    assign layer_1_weights[29][67] = 6'sd6;
    assign layer_1_weights[29][68] = 6'sd3;
    assign layer_1_weights[29][69] = 6'sd2;
    assign layer_1_weights[29][70] = -6'sd1;
    assign layer_1_weights[29][71] = -6'sd4;
    assign layer_1_weights[29][72] = 6'sd0;
    assign layer_1_weights[29][73] = -6'sd4;
    assign layer_1_weights[29][74] = 6'sd1;
    assign layer_1_weights[29][75] = -6'sd1;
    assign layer_1_weights[29][76] = -6'sd1;
    assign layer_1_weights[29][77] = -6'sd2;
    assign layer_1_weights[29][78] = 6'sd2;
    assign layer_1_weights[29][79] = 6'sd3;
    assign layer_1_weights[29][80] = 6'sd6;
    assign layer_1_weights[29][81] = 6'sd4;
    assign layer_1_weights[29][82] = 6'sd4;
    assign layer_1_weights[29][83] = 6'sd1;
    assign layer_1_weights[29][84] = 6'sd3;
    assign layer_1_weights[29][85] = 6'sd4;
    assign layer_1_weights[29][86] = 6'sd4;
    assign layer_1_weights[29][87] = 6'sd1;
    assign layer_1_weights[29][88] = 6'sd1;
    assign layer_1_weights[29][89] = -6'sd3;
    assign layer_1_weights[29][90] = -6'sd1;
    assign layer_1_weights[29][91] = 6'sd3;
    assign layer_1_weights[29][92] = 6'sd3;
    assign layer_1_weights[29][93] = -6'sd1;
    assign layer_1_weights[29][94] = -6'sd1;
    assign layer_1_weights[29][95] = 6'sd3;
    assign layer_1_weights[29][96] = -6'sd1;
    assign layer_1_weights[29][97] = 6'sd3;
    assign layer_1_weights[29][98] = 6'sd2;
    assign layer_1_weights[29][99] = 6'sd2;
    assign layer_1_weights[29][100] = 6'sd2;
    assign layer_1_weights[29][101] = 6'sd5;
    assign layer_1_weights[29][102] = 6'sd7;
    assign layer_1_weights[29][103] = 6'sd1;
    assign layer_1_weights[29][104] = -6'sd5;
    assign layer_1_weights[29][105] = -6'sd2;
    assign layer_1_weights[29][106] = -6'sd5;
    assign layer_1_weights[29][107] = -6'sd2;
    assign layer_1_weights[29][108] = 6'sd4;
    assign layer_1_weights[29][109] = -6'sd7;
    assign layer_1_weights[29][110] = -6'sd2;
    assign layer_1_weights[29][111] = 6'sd2;
    assign layer_1_weights[29][112] = 6'sd2;
    assign layer_1_weights[29][113] = 6'sd4;
    assign layer_1_weights[29][114] = -6'sd3;
    assign layer_1_weights[29][115] = -6'sd3;
    assign layer_1_weights[29][116] = -6'sd4;
    assign layer_1_weights[29][117] = -6'sd5;
    assign layer_1_weights[29][118] = -6'sd9;
    assign layer_1_weights[29][119] = 6'sd1;
    assign layer_1_weights[29][120] = 6'sd0;
    assign layer_1_weights[29][121] = -6'sd9;
    assign layer_1_weights[29][122] = -6'sd6;
    assign layer_1_weights[29][123] = -6'sd9;
    assign layer_1_weights[29][124] = -6'sd8;
    assign layer_1_weights[29][125] = -6'sd11;
    assign layer_1_weights[29][126] = -6'sd14;
    assign layer_1_weights[29][127] = -6'sd17;
    assign layer_1_weights[29][128] = -6'sd14;
    assign layer_1_weights[29][129] = -6'sd3;
    assign layer_1_weights[29][130] = -6'sd9;
    assign layer_1_weights[29][131] = 6'sd1;
    assign layer_1_weights[29][132] = 6'sd1;
    assign layer_1_weights[29][133] = -6'sd2;
    assign layer_1_weights[29][134] = -6'sd8;
    assign layer_1_weights[29][135] = -6'sd11;
    assign layer_1_weights[29][136] = -6'sd6;
    assign layer_1_weights[29][137] = -6'sd14;
    assign layer_1_weights[29][138] = -6'sd7;
    assign layer_1_weights[29][139] = 6'sd3;
    assign layer_1_weights[29][140] = -6'sd6;
    assign layer_1_weights[29][141] = -6'sd6;
    assign layer_1_weights[29][142] = 6'sd0;
    assign layer_1_weights[29][143] = 6'sd0;
    assign layer_1_biases[29] = 6'sd0;
    assign layer_1_weights[30][0] = -6'sd1;
    assign layer_1_weights[30][1] = -6'sd2;
    assign layer_1_weights[30][2] = 6'sd3;
    assign layer_1_weights[30][3] = 6'sd5;
    assign layer_1_weights[30][4] = 6'sd3;
    assign layer_1_weights[30][5] = 6'sd4;
    assign layer_1_weights[30][6] = -6'sd1;
    assign layer_1_weights[30][7] = 6'sd7;
    assign layer_1_weights[30][8] = 6'sd2;
    assign layer_1_weights[30][9] = 6'sd9;
    assign layer_1_weights[30][10] = -6'sd1;
    assign layer_1_weights[30][11] = -6'sd1;
    assign layer_1_weights[30][12] = -6'sd2;
    assign layer_1_weights[30][13] = 6'sd1;
    assign layer_1_weights[30][14] = 6'sd7;
    assign layer_1_weights[30][15] = 6'sd5;
    assign layer_1_weights[30][16] = 6'sd2;
    assign layer_1_weights[30][17] = 6'sd1;
    assign layer_1_weights[30][18] = -6'sd2;
    assign layer_1_weights[30][19] = 6'sd0;
    assign layer_1_weights[30][20] = -6'sd4;
    assign layer_1_weights[30][21] = -6'sd3;
    assign layer_1_weights[30][22] = -6'sd2;
    assign layer_1_weights[30][23] = 6'sd0;
    assign layer_1_weights[30][24] = -6'sd1;
    assign layer_1_weights[30][25] = 6'sd2;
    assign layer_1_weights[30][26] = 6'sd2;
    assign layer_1_weights[30][27] = 6'sd0;
    assign layer_1_weights[30][28] = -6'sd1;
    assign layer_1_weights[30][29] = 6'sd1;
    assign layer_1_weights[30][30] = -6'sd1;
    assign layer_1_weights[30][31] = 6'sd0;
    assign layer_1_weights[30][32] = -6'sd1;
    assign layer_1_weights[30][33] = -6'sd7;
    assign layer_1_weights[30][34] = -6'sd3;
    assign layer_1_weights[30][35] = -6'sd3;
    assign layer_1_weights[30][36] = -6'sd2;
    assign layer_1_weights[30][37] = 6'sd12;
    assign layer_1_weights[30][38] = 6'sd3;
    assign layer_1_weights[30][39] = -6'sd1;
    assign layer_1_weights[30][40] = 6'sd0;
    assign layer_1_weights[30][41] = 6'sd1;
    assign layer_1_weights[30][42] = 6'sd6;
    assign layer_1_weights[30][43] = 6'sd6;
    assign layer_1_weights[30][44] = 6'sd6;
    assign layer_1_weights[30][45] = 6'sd2;
    assign layer_1_weights[30][46] = -6'sd3;
    assign layer_1_weights[30][47] = -6'sd5;
    assign layer_1_weights[30][48] = -6'sd2;
    assign layer_1_weights[30][49] = 6'sd0;
    assign layer_1_weights[30][50] = 6'sd2;
    assign layer_1_weights[30][51] = -6'sd2;
    assign layer_1_weights[30][52] = -6'sd3;
    assign layer_1_weights[30][53] = 6'sd1;
    assign layer_1_weights[30][54] = -6'sd2;
    assign layer_1_weights[30][55] = 6'sd1;
    assign layer_1_weights[30][56] = 6'sd7;
    assign layer_1_weights[30][57] = 6'sd5;
    assign layer_1_weights[30][58] = -6'sd4;
    assign layer_1_weights[30][59] = -6'sd11;
    assign layer_1_weights[30][60] = -6'sd11;
    assign layer_1_weights[30][61] = 6'sd2;
    assign layer_1_weights[30][62] = 6'sd0;
    assign layer_1_weights[30][63] = 6'sd1;
    assign layer_1_weights[30][64] = 6'sd0;
    assign layer_1_weights[30][65] = -6'sd1;
    assign layer_1_weights[30][66] = -6'sd5;
    assign layer_1_weights[30][67] = -6'sd2;
    assign layer_1_weights[30][68] = 6'sd1;
    assign layer_1_weights[30][69] = 6'sd2;
    assign layer_1_weights[30][70] = -6'sd2;
    assign layer_1_weights[30][71] = -6'sd12;
    assign layer_1_weights[30][72] = 6'sd2;
    assign layer_1_weights[30][73] = -6'sd2;
    assign layer_1_weights[30][74] = -6'sd3;
    assign layer_1_weights[30][75] = -6'sd3;
    assign layer_1_weights[30][76] = 6'sd3;
    assign layer_1_weights[30][77] = 6'sd4;
    assign layer_1_weights[30][78] = -6'sd2;
    assign layer_1_weights[30][79] = 6'sd0;
    assign layer_1_weights[30][80] = 6'sd3;
    assign layer_1_weights[30][81] = 6'sd2;
    assign layer_1_weights[30][82] = 6'sd5;
    assign layer_1_weights[30][83] = -6'sd5;
    assign layer_1_weights[30][84] = 6'sd6;
    assign layer_1_weights[30][85] = 6'sd0;
    assign layer_1_weights[30][86] = -6'sd1;
    assign layer_1_weights[30][87] = 6'sd1;
    assign layer_1_weights[30][88] = 6'sd1;
    assign layer_1_weights[30][89] = 6'sd6;
    assign layer_1_weights[30][90] = 6'sd1;
    assign layer_1_weights[30][91] = 6'sd0;
    assign layer_1_weights[30][92] = 6'sd2;
    assign layer_1_weights[30][93] = -6'sd2;
    assign layer_1_weights[30][94] = 6'sd0;
    assign layer_1_weights[30][95] = -6'sd1;
    assign layer_1_weights[30][96] = 6'sd7;
    assign layer_1_weights[30][97] = -6'sd2;
    assign layer_1_weights[30][98] = -6'sd3;
    assign layer_1_weights[30][99] = -6'sd1;
    assign layer_1_weights[30][100] = 6'sd3;
    assign layer_1_weights[30][101] = 6'sd4;
    assign layer_1_weights[30][102] = 6'sd0;
    assign layer_1_weights[30][103] = 6'sd2;
    assign layer_1_weights[30][104] = 6'sd2;
    assign layer_1_weights[30][105] = 6'sd1;
    assign layer_1_weights[30][106] = -6'sd7;
    assign layer_1_weights[30][107] = -6'sd2;
    assign layer_1_weights[30][108] = 6'sd1;
    assign layer_1_weights[30][109] = -6'sd2;
    assign layer_1_weights[30][110] = -6'sd2;
    assign layer_1_weights[30][111] = -6'sd2;
    assign layer_1_weights[30][112] = 6'sd1;
    assign layer_1_weights[30][113] = 6'sd3;
    assign layer_1_weights[30][114] = 6'sd1;
    assign layer_1_weights[30][115] = 6'sd2;
    assign layer_1_weights[30][116] = 6'sd3;
    assign layer_1_weights[30][117] = -6'sd4;
    assign layer_1_weights[30][118] = -6'sd1;
    assign layer_1_weights[30][119] = -6'sd6;
    assign layer_1_weights[30][120] = 6'sd1;
    assign layer_1_weights[30][121] = 6'sd8;
    assign layer_1_weights[30][122] = 6'sd0;
    assign layer_1_weights[30][123] = 6'sd1;
    assign layer_1_weights[30][124] = 6'sd3;
    assign layer_1_weights[30][125] = 6'sd2;
    assign layer_1_weights[30][126] = 6'sd0;
    assign layer_1_weights[30][127] = -6'sd1;
    assign layer_1_weights[30][128] = 6'sd2;
    assign layer_1_weights[30][129] = 6'sd3;
    assign layer_1_weights[30][130] = -6'sd3;
    assign layer_1_weights[30][131] = 6'sd4;
    assign layer_1_weights[30][132] = 6'sd1;
    assign layer_1_weights[30][133] = 6'sd5;
    assign layer_1_weights[30][134] = 6'sd5;
    assign layer_1_weights[30][135] = 6'sd7;
    assign layer_1_weights[30][136] = 6'sd6;
    assign layer_1_weights[30][137] = 6'sd4;
    assign layer_1_weights[30][138] = -6'sd3;
    assign layer_1_weights[30][139] = 6'sd0;
    assign layer_1_weights[30][140] = -6'sd1;
    assign layer_1_weights[30][141] = -6'sd1;
    assign layer_1_weights[30][142] = -6'sd1;
    assign layer_1_weights[30][143] = -6'sd1;
    assign layer_1_biases[30] = -6'sd4;
    assign layer_1_weights[31][0] = 6'sd1;
    assign layer_1_weights[31][1] = 6'sd2;
    assign layer_1_weights[31][2] = 6'sd0;
    assign layer_1_weights[31][3] = -6'sd1;
    assign layer_1_weights[31][4] = -6'sd7;
    assign layer_1_weights[31][5] = -6'sd2;
    assign layer_1_weights[31][6] = 6'sd0;
    assign layer_1_weights[31][7] = -6'sd3;
    assign layer_1_weights[31][8] = -6'sd11;
    assign layer_1_weights[31][9] = -6'sd9;
    assign layer_1_weights[31][10] = -6'sd2;
    assign layer_1_weights[31][11] = 6'sd0;
    assign layer_1_weights[31][12] = 6'sd0;
    assign layer_1_weights[31][13] = -6'sd1;
    assign layer_1_weights[31][14] = -6'sd6;
    assign layer_1_weights[31][15] = -6'sd16;
    assign layer_1_weights[31][16] = -6'sd11;
    assign layer_1_weights[31][17] = -6'sd3;
    assign layer_1_weights[31][18] = -6'sd3;
    assign layer_1_weights[31][19] = 6'sd0;
    assign layer_1_weights[31][20] = -6'sd2;
    assign layer_1_weights[31][21] = -6'sd4;
    assign layer_1_weights[31][22] = -6'sd4;
    assign layer_1_weights[31][23] = -6'sd5;
    assign layer_1_weights[31][24] = 6'sd0;
    assign layer_1_weights[31][25] = -6'sd6;
    assign layer_1_weights[31][26] = 6'sd1;
    assign layer_1_weights[31][27] = -6'sd2;
    assign layer_1_weights[31][28] = 6'sd1;
    assign layer_1_weights[31][29] = 6'sd2;
    assign layer_1_weights[31][30] = -6'sd2;
    assign layer_1_weights[31][31] = 6'sd0;
    assign layer_1_weights[31][32] = 6'sd3;
    assign layer_1_weights[31][33] = 6'sd0;
    assign layer_1_weights[31][34] = -6'sd1;
    assign layer_1_weights[31][35] = -6'sd3;
    assign layer_1_weights[31][36] = 6'sd2;
    assign layer_1_weights[31][37] = -6'sd2;
    assign layer_1_weights[31][38] = -6'sd2;
    assign layer_1_weights[31][39] = 6'sd2;
    assign layer_1_weights[31][40] = 6'sd1;
    assign layer_1_weights[31][41] = 6'sd0;
    assign layer_1_weights[31][42] = -6'sd2;
    assign layer_1_weights[31][43] = 6'sd4;
    assign layer_1_weights[31][44] = 6'sd5;
    assign layer_1_weights[31][45] = 6'sd4;
    assign layer_1_weights[31][46] = 6'sd0;
    assign layer_1_weights[31][47] = 6'sd2;
    assign layer_1_weights[31][48] = 6'sd0;
    assign layer_1_weights[31][49] = 6'sd1;
    assign layer_1_weights[31][50] = 6'sd2;
    assign layer_1_weights[31][51] = 6'sd2;
    assign layer_1_weights[31][52] = -6'sd3;
    assign layer_1_weights[31][53] = -6'sd3;
    assign layer_1_weights[31][54] = 6'sd0;
    assign layer_1_weights[31][55] = 6'sd7;
    assign layer_1_weights[31][56] = 6'sd6;
    assign layer_1_weights[31][57] = -6'sd1;
    assign layer_1_weights[31][58] = -6'sd4;
    assign layer_1_weights[31][59] = 6'sd0;
    assign layer_1_weights[31][60] = 6'sd4;
    assign layer_1_weights[31][61] = -6'sd6;
    assign layer_1_weights[31][62] = -6'sd1;
    assign layer_1_weights[31][63] = -6'sd1;
    assign layer_1_weights[31][64] = 6'sd2;
    assign layer_1_weights[31][65] = 6'sd2;
    assign layer_1_weights[31][66] = 6'sd0;
    assign layer_1_weights[31][67] = 6'sd8;
    assign layer_1_weights[31][68] = 6'sd3;
    assign layer_1_weights[31][69] = 6'sd1;
    assign layer_1_weights[31][70] = -6'sd3;
    assign layer_1_weights[31][71] = -6'sd1;
    assign layer_1_weights[31][72] = 6'sd5;
    assign layer_1_weights[31][73] = 6'sd1;
    assign layer_1_weights[31][74] = 6'sd0;
    assign layer_1_weights[31][75] = -6'sd1;
    assign layer_1_weights[31][76] = 6'sd1;
    assign layer_1_weights[31][77] = 6'sd1;
    assign layer_1_weights[31][78] = 6'sd3;
    assign layer_1_weights[31][79] = 6'sd5;
    assign layer_1_weights[31][80] = 6'sd1;
    assign layer_1_weights[31][81] = -6'sd1;
    assign layer_1_weights[31][82] = -6'sd2;
    assign layer_1_weights[31][83] = -6'sd7;
    assign layer_1_weights[31][84] = 6'sd6;
    assign layer_1_weights[31][85] = -6'sd1;
    assign layer_1_weights[31][86] = -6'sd2;
    assign layer_1_weights[31][87] = -6'sd1;
    assign layer_1_weights[31][88] = 6'sd1;
    assign layer_1_weights[31][89] = 6'sd4;
    assign layer_1_weights[31][90] = 6'sd0;
    assign layer_1_weights[31][91] = 6'sd0;
    assign layer_1_weights[31][92] = -6'sd5;
    assign layer_1_weights[31][93] = -6'sd6;
    assign layer_1_weights[31][94] = -6'sd6;
    assign layer_1_weights[31][95] = 6'sd1;
    assign layer_1_weights[31][96] = 6'sd4;
    assign layer_1_weights[31][97] = 6'sd0;
    assign layer_1_weights[31][98] = -6'sd4;
    assign layer_1_weights[31][99] = -6'sd3;
    assign layer_1_weights[31][100] = 6'sd0;
    assign layer_1_weights[31][101] = 6'sd3;
    assign layer_1_weights[31][102] = -6'sd3;
    assign layer_1_weights[31][103] = -6'sd7;
    assign layer_1_weights[31][104] = -6'sd3;
    assign layer_1_weights[31][105] = -6'sd8;
    assign layer_1_weights[31][106] = -6'sd10;
    assign layer_1_weights[31][107] = 6'sd5;
    assign layer_1_weights[31][108] = 6'sd0;
    assign layer_1_weights[31][109] = -6'sd7;
    assign layer_1_weights[31][110] = -6'sd2;
    assign layer_1_weights[31][111] = -6'sd4;
    assign layer_1_weights[31][112] = 6'sd3;
    assign layer_1_weights[31][113] = 6'sd6;
    assign layer_1_weights[31][114] = -6'sd6;
    assign layer_1_weights[31][115] = -6'sd9;
    assign layer_1_weights[31][116] = -6'sd12;
    assign layer_1_weights[31][117] = 6'sd0;
    assign layer_1_weights[31][118] = -6'sd1;
    assign layer_1_weights[31][119] = 6'sd5;
    assign layer_1_weights[31][120] = -6'sd2;
    assign layer_1_weights[31][121] = 6'sd2;
    assign layer_1_weights[31][122] = 6'sd1;
    assign layer_1_weights[31][123] = -6'sd1;
    assign layer_1_weights[31][124] = 6'sd2;
    assign layer_1_weights[31][125] = 6'sd2;
    assign layer_1_weights[31][126] = 6'sd0;
    assign layer_1_weights[31][127] = -6'sd14;
    assign layer_1_weights[31][128] = -6'sd16;
    assign layer_1_weights[31][129] = 6'sd0;
    assign layer_1_weights[31][130] = 6'sd1;
    assign layer_1_weights[31][131] = -6'sd1;
    assign layer_1_weights[31][132] = -6'sd1;
    assign layer_1_weights[31][133] = 6'sd1;
    assign layer_1_weights[31][134] = 6'sd1;
    assign layer_1_weights[31][135] = 6'sd1;
    assign layer_1_weights[31][136] = -6'sd2;
    assign layer_1_weights[31][137] = 6'sd0;
    assign layer_1_weights[31][138] = -6'sd5;
    assign layer_1_weights[31][139] = -6'sd2;
    assign layer_1_weights[31][140] = -6'sd8;
    assign layer_1_weights[31][141] = -6'sd7;
    assign layer_1_weights[31][142] = 6'sd0;
    assign layer_1_weights[31][143] = 6'sd1;
    assign layer_1_biases[31] = -6'sd2;

    wire signed [5:0] layer_1_output_0;
    wire signed [5:0] layer_1_output_1;
    wire signed [5:0] layer_1_output_2;
    wire signed [5:0] layer_1_output_3;
    wire signed [5:0] layer_1_output_4;
    wire signed [5:0] layer_1_output_5;
    wire signed [5:0] layer_1_output_6;
    wire signed [5:0] layer_1_output_7;
    wire signed [5:0] layer_1_output_8;
    wire signed [5:0] layer_1_output_9;
    wire signed [5:0] layer_1_output_10;
    wire signed [5:0] layer_1_output_11;
    wire signed [5:0] layer_1_output_12;
    wire signed [5:0] layer_1_output_13;
    wire signed [5:0] layer_1_output_14;
    wire signed [5:0] layer_1_output_15;
    wire signed [5:0] layer_1_output_16;
    wire signed [5:0] layer_1_output_17;
    wire signed [5:0] layer_1_output_18;
    wire signed [5:0] layer_1_output_19;
    wire signed [5:0] layer_1_output_20;
    wire signed [5:0] layer_1_output_21;
    wire signed [5:0] layer_1_output_22;
    wire signed [5:0] layer_1_output_23;
    wire signed [5:0] layer_1_output_24;
    wire signed [5:0] layer_1_output_25;
    wire signed [5:0] layer_1_output_26;
    wire signed [5:0] layer_1_output_27;
    wire signed [5:0] layer_1_output_28;
    wire signed [5:0] layer_1_output_29;
    wire signed [5:0] layer_1_output_30;
    wire signed [5:0] layer_1_output_31;
    assign layer_1_output_0 = relu(layer_1_biases[0] + inp[0] * layer_1_weights[0][0] + inp[1] * layer_1_weights[0][1] + inp[2] * layer_1_weights[0][2] + inp[3] * layer_1_weights[0][3] + inp[4] * layer_1_weights[0][4] + inp[5] * layer_1_weights[0][5] + inp[6] * layer_1_weights[0][6] + inp[7] * layer_1_weights[0][7] + inp[8] * layer_1_weights[0][8] + inp[9] * layer_1_weights[0][9] + inp[10] * layer_1_weights[0][10] + inp[11] * layer_1_weights[0][11] + inp[12] * layer_1_weights[0][12] + inp[13] * layer_1_weights[0][13] + inp[14] * layer_1_weights[0][14] + inp[15] * layer_1_weights[0][15] + inp[16] * layer_1_weights[0][16] + inp[17] * layer_1_weights[0][17] + inp[18] * layer_1_weights[0][18] + inp[19] * layer_1_weights[0][19] + inp[20] * layer_1_weights[0][20] + inp[21] * layer_1_weights[0][21] + inp[22] * layer_1_weights[0][22] + inp[23] * layer_1_weights[0][23] + inp[24] * layer_1_weights[0][24] + inp[25] * layer_1_weights[0][25] + inp[26] * layer_1_weights[0][26] + inp[27] * layer_1_weights[0][27] + inp[28] * layer_1_weights[0][28] + inp[29] * layer_1_weights[0][29] + inp[30] * layer_1_weights[0][30] + inp[31] * layer_1_weights[0][31] + inp[32] * layer_1_weights[0][32] + inp[33] * layer_1_weights[0][33] + inp[34] * layer_1_weights[0][34] + inp[35] * layer_1_weights[0][35] + inp[36] * layer_1_weights[0][36] + inp[37] * layer_1_weights[0][37] + inp[38] * layer_1_weights[0][38] + inp[39] * layer_1_weights[0][39] + inp[40] * layer_1_weights[0][40] + inp[41] * layer_1_weights[0][41] + inp[42] * layer_1_weights[0][42] + inp[43] * layer_1_weights[0][43] + inp[44] * layer_1_weights[0][44] + inp[45] * layer_1_weights[0][45] + inp[46] * layer_1_weights[0][46] + inp[47] * layer_1_weights[0][47] + inp[48] * layer_1_weights[0][48] + inp[49] * layer_1_weights[0][49] + inp[50] * layer_1_weights[0][50] + inp[51] * layer_1_weights[0][51] + inp[52] * layer_1_weights[0][52] + inp[53] * layer_1_weights[0][53] + inp[54] * layer_1_weights[0][54] + inp[55] * layer_1_weights[0][55] + inp[56] * layer_1_weights[0][56] + inp[57] * layer_1_weights[0][57] + inp[58] * layer_1_weights[0][58] + inp[59] * layer_1_weights[0][59] + inp[60] * layer_1_weights[0][60] + inp[61] * layer_1_weights[0][61] + inp[62] * layer_1_weights[0][62] + inp[63] * layer_1_weights[0][63] + inp[64] * layer_1_weights[0][64] + inp[65] * layer_1_weights[0][65] + inp[66] * layer_1_weights[0][66] + inp[67] * layer_1_weights[0][67] + inp[68] * layer_1_weights[0][68] + inp[69] * layer_1_weights[0][69] + inp[70] * layer_1_weights[0][70] + inp[71] * layer_1_weights[0][71] + inp[72] * layer_1_weights[0][72] + inp[73] * layer_1_weights[0][73] + inp[74] * layer_1_weights[0][74] + inp[75] * layer_1_weights[0][75] + inp[76] * layer_1_weights[0][76] + inp[77] * layer_1_weights[0][77] + inp[78] * layer_1_weights[0][78] + inp[79] * layer_1_weights[0][79] + inp[80] * layer_1_weights[0][80] + inp[81] * layer_1_weights[0][81] + inp[82] * layer_1_weights[0][82] + inp[83] * layer_1_weights[0][83] + inp[84] * layer_1_weights[0][84] + inp[85] * layer_1_weights[0][85] + inp[86] * layer_1_weights[0][86] + inp[87] * layer_1_weights[0][87] + inp[88] * layer_1_weights[0][88] + inp[89] * layer_1_weights[0][89] + inp[90] * layer_1_weights[0][90] + inp[91] * layer_1_weights[0][91] + inp[92] * layer_1_weights[0][92] + inp[93] * layer_1_weights[0][93] + inp[94] * layer_1_weights[0][94] + inp[95] * layer_1_weights[0][95] + inp[96] * layer_1_weights[0][96] + inp[97] * layer_1_weights[0][97] + inp[98] * layer_1_weights[0][98] + inp[99] * layer_1_weights[0][99] + inp[100] * layer_1_weights[0][100] + inp[101] * layer_1_weights[0][101] + inp[102] * layer_1_weights[0][102] + inp[103] * layer_1_weights[0][103] + inp[104] * layer_1_weights[0][104] + inp[105] * layer_1_weights[0][105] + inp[106] * layer_1_weights[0][106] + inp[107] * layer_1_weights[0][107] + inp[108] * layer_1_weights[0][108] + inp[109] * layer_1_weights[0][109] + inp[110] * layer_1_weights[0][110] + inp[111] * layer_1_weights[0][111] + inp[112] * layer_1_weights[0][112] + inp[113] * layer_1_weights[0][113] + inp[114] * layer_1_weights[0][114] + inp[115] * layer_1_weights[0][115] + inp[116] * layer_1_weights[0][116] + inp[117] * layer_1_weights[0][117] + inp[118] * layer_1_weights[0][118] + inp[119] * layer_1_weights[0][119] + inp[120] * layer_1_weights[0][120] + inp[121] * layer_1_weights[0][121] + inp[122] * layer_1_weights[0][122] + inp[123] * layer_1_weights[0][123] + inp[124] * layer_1_weights[0][124] + inp[125] * layer_1_weights[0][125] + inp[126] * layer_1_weights[0][126] + inp[127] * layer_1_weights[0][127] + inp[128] * layer_1_weights[0][128] + inp[129] * layer_1_weights[0][129] + inp[130] * layer_1_weights[0][130] + inp[131] * layer_1_weights[0][131] + inp[132] * layer_1_weights[0][132] + inp[133] * layer_1_weights[0][133] + inp[134] * layer_1_weights[0][134] + inp[135] * layer_1_weights[0][135] + inp[136] * layer_1_weights[0][136] + inp[137] * layer_1_weights[0][137] + inp[138] * layer_1_weights[0][138] + inp[139] * layer_1_weights[0][139] + inp[140] * layer_1_weights[0][140] + inp[141] * layer_1_weights[0][141] + inp[142] * layer_1_weights[0][142] + inp[143] * layer_1_weights[0][143]);
    assign layer_1_output_1 = relu(layer_1_biases[1] + inp[0] * layer_1_weights[1][0] + inp[1] * layer_1_weights[1][1] + inp[2] * layer_1_weights[1][2] + inp[3] * layer_1_weights[1][3] + inp[4] * layer_1_weights[1][4] + inp[5] * layer_1_weights[1][5] + inp[6] * layer_1_weights[1][6] + inp[7] * layer_1_weights[1][7] + inp[8] * layer_1_weights[1][8] + inp[9] * layer_1_weights[1][9] + inp[10] * layer_1_weights[1][10] + inp[11] * layer_1_weights[1][11] + inp[12] * layer_1_weights[1][12] + inp[13] * layer_1_weights[1][13] + inp[14] * layer_1_weights[1][14] + inp[15] * layer_1_weights[1][15] + inp[16] * layer_1_weights[1][16] + inp[17] * layer_1_weights[1][17] + inp[18] * layer_1_weights[1][18] + inp[19] * layer_1_weights[1][19] + inp[20] * layer_1_weights[1][20] + inp[21] * layer_1_weights[1][21] + inp[22] * layer_1_weights[1][22] + inp[23] * layer_1_weights[1][23] + inp[24] * layer_1_weights[1][24] + inp[25] * layer_1_weights[1][25] + inp[26] * layer_1_weights[1][26] + inp[27] * layer_1_weights[1][27] + inp[28] * layer_1_weights[1][28] + inp[29] * layer_1_weights[1][29] + inp[30] * layer_1_weights[1][30] + inp[31] * layer_1_weights[1][31] + inp[32] * layer_1_weights[1][32] + inp[33] * layer_1_weights[1][33] + inp[34] * layer_1_weights[1][34] + inp[35] * layer_1_weights[1][35] + inp[36] * layer_1_weights[1][36] + inp[37] * layer_1_weights[1][37] + inp[38] * layer_1_weights[1][38] + inp[39] * layer_1_weights[1][39] + inp[40] * layer_1_weights[1][40] + inp[41] * layer_1_weights[1][41] + inp[42] * layer_1_weights[1][42] + inp[43] * layer_1_weights[1][43] + inp[44] * layer_1_weights[1][44] + inp[45] * layer_1_weights[1][45] + inp[46] * layer_1_weights[1][46] + inp[47] * layer_1_weights[1][47] + inp[48] * layer_1_weights[1][48] + inp[49] * layer_1_weights[1][49] + inp[50] * layer_1_weights[1][50] + inp[51] * layer_1_weights[1][51] + inp[52] * layer_1_weights[1][52] + inp[53] * layer_1_weights[1][53] + inp[54] * layer_1_weights[1][54] + inp[55] * layer_1_weights[1][55] + inp[56] * layer_1_weights[1][56] + inp[57] * layer_1_weights[1][57] + inp[58] * layer_1_weights[1][58] + inp[59] * layer_1_weights[1][59] + inp[60] * layer_1_weights[1][60] + inp[61] * layer_1_weights[1][61] + inp[62] * layer_1_weights[1][62] + inp[63] * layer_1_weights[1][63] + inp[64] * layer_1_weights[1][64] + inp[65] * layer_1_weights[1][65] + inp[66] * layer_1_weights[1][66] + inp[67] * layer_1_weights[1][67] + inp[68] * layer_1_weights[1][68] + inp[69] * layer_1_weights[1][69] + inp[70] * layer_1_weights[1][70] + inp[71] * layer_1_weights[1][71] + inp[72] * layer_1_weights[1][72] + inp[73] * layer_1_weights[1][73] + inp[74] * layer_1_weights[1][74] + inp[75] * layer_1_weights[1][75] + inp[76] * layer_1_weights[1][76] + inp[77] * layer_1_weights[1][77] + inp[78] * layer_1_weights[1][78] + inp[79] * layer_1_weights[1][79] + inp[80] * layer_1_weights[1][80] + inp[81] * layer_1_weights[1][81] + inp[82] * layer_1_weights[1][82] + inp[83] * layer_1_weights[1][83] + inp[84] * layer_1_weights[1][84] + inp[85] * layer_1_weights[1][85] + inp[86] * layer_1_weights[1][86] + inp[87] * layer_1_weights[1][87] + inp[88] * layer_1_weights[1][88] + inp[89] * layer_1_weights[1][89] + inp[90] * layer_1_weights[1][90] + inp[91] * layer_1_weights[1][91] + inp[92] * layer_1_weights[1][92] + inp[93] * layer_1_weights[1][93] + inp[94] * layer_1_weights[1][94] + inp[95] * layer_1_weights[1][95] + inp[96] * layer_1_weights[1][96] + inp[97] * layer_1_weights[1][97] + inp[98] * layer_1_weights[1][98] + inp[99] * layer_1_weights[1][99] + inp[100] * layer_1_weights[1][100] + inp[101] * layer_1_weights[1][101] + inp[102] * layer_1_weights[1][102] + inp[103] * layer_1_weights[1][103] + inp[104] * layer_1_weights[1][104] + inp[105] * layer_1_weights[1][105] + inp[106] * layer_1_weights[1][106] + inp[107] * layer_1_weights[1][107] + inp[108] * layer_1_weights[1][108] + inp[109] * layer_1_weights[1][109] + inp[110] * layer_1_weights[1][110] + inp[111] * layer_1_weights[1][111] + inp[112] * layer_1_weights[1][112] + inp[113] * layer_1_weights[1][113] + inp[114] * layer_1_weights[1][114] + inp[115] * layer_1_weights[1][115] + inp[116] * layer_1_weights[1][116] + inp[117] * layer_1_weights[1][117] + inp[118] * layer_1_weights[1][118] + inp[119] * layer_1_weights[1][119] + inp[120] * layer_1_weights[1][120] + inp[121] * layer_1_weights[1][121] + inp[122] * layer_1_weights[1][122] + inp[123] * layer_1_weights[1][123] + inp[124] * layer_1_weights[1][124] + inp[125] * layer_1_weights[1][125] + inp[126] * layer_1_weights[1][126] + inp[127] * layer_1_weights[1][127] + inp[128] * layer_1_weights[1][128] + inp[129] * layer_1_weights[1][129] + inp[130] * layer_1_weights[1][130] + inp[131] * layer_1_weights[1][131] + inp[132] * layer_1_weights[1][132] + inp[133] * layer_1_weights[1][133] + inp[134] * layer_1_weights[1][134] + inp[135] * layer_1_weights[1][135] + inp[136] * layer_1_weights[1][136] + inp[137] * layer_1_weights[1][137] + inp[138] * layer_1_weights[1][138] + inp[139] * layer_1_weights[1][139] + inp[140] * layer_1_weights[1][140] + inp[141] * layer_1_weights[1][141] + inp[142] * layer_1_weights[1][142] + inp[143] * layer_1_weights[1][143]);
    assign layer_1_output_2 = relu(layer_1_biases[2] + inp[0] * layer_1_weights[2][0] + inp[1] * layer_1_weights[2][1] + inp[2] * layer_1_weights[2][2] + inp[3] * layer_1_weights[2][3] + inp[4] * layer_1_weights[2][4] + inp[5] * layer_1_weights[2][5] + inp[6] * layer_1_weights[2][6] + inp[7] * layer_1_weights[2][7] + inp[8] * layer_1_weights[2][8] + inp[9] * layer_1_weights[2][9] + inp[10] * layer_1_weights[2][10] + inp[11] * layer_1_weights[2][11] + inp[12] * layer_1_weights[2][12] + inp[13] * layer_1_weights[2][13] + inp[14] * layer_1_weights[2][14] + inp[15] * layer_1_weights[2][15] + inp[16] * layer_1_weights[2][16] + inp[17] * layer_1_weights[2][17] + inp[18] * layer_1_weights[2][18] + inp[19] * layer_1_weights[2][19] + inp[20] * layer_1_weights[2][20] + inp[21] * layer_1_weights[2][21] + inp[22] * layer_1_weights[2][22] + inp[23] * layer_1_weights[2][23] + inp[24] * layer_1_weights[2][24] + inp[25] * layer_1_weights[2][25] + inp[26] * layer_1_weights[2][26] + inp[27] * layer_1_weights[2][27] + inp[28] * layer_1_weights[2][28] + inp[29] * layer_1_weights[2][29] + inp[30] * layer_1_weights[2][30] + inp[31] * layer_1_weights[2][31] + inp[32] * layer_1_weights[2][32] + inp[33] * layer_1_weights[2][33] + inp[34] * layer_1_weights[2][34] + inp[35] * layer_1_weights[2][35] + inp[36] * layer_1_weights[2][36] + inp[37] * layer_1_weights[2][37] + inp[38] * layer_1_weights[2][38] + inp[39] * layer_1_weights[2][39] + inp[40] * layer_1_weights[2][40] + inp[41] * layer_1_weights[2][41] + inp[42] * layer_1_weights[2][42] + inp[43] * layer_1_weights[2][43] + inp[44] * layer_1_weights[2][44] + inp[45] * layer_1_weights[2][45] + inp[46] * layer_1_weights[2][46] + inp[47] * layer_1_weights[2][47] + inp[48] * layer_1_weights[2][48] + inp[49] * layer_1_weights[2][49] + inp[50] * layer_1_weights[2][50] + inp[51] * layer_1_weights[2][51] + inp[52] * layer_1_weights[2][52] + inp[53] * layer_1_weights[2][53] + inp[54] * layer_1_weights[2][54] + inp[55] * layer_1_weights[2][55] + inp[56] * layer_1_weights[2][56] + inp[57] * layer_1_weights[2][57] + inp[58] * layer_1_weights[2][58] + inp[59] * layer_1_weights[2][59] + inp[60] * layer_1_weights[2][60] + inp[61] * layer_1_weights[2][61] + inp[62] * layer_1_weights[2][62] + inp[63] * layer_1_weights[2][63] + inp[64] * layer_1_weights[2][64] + inp[65] * layer_1_weights[2][65] + inp[66] * layer_1_weights[2][66] + inp[67] * layer_1_weights[2][67] + inp[68] * layer_1_weights[2][68] + inp[69] * layer_1_weights[2][69] + inp[70] * layer_1_weights[2][70] + inp[71] * layer_1_weights[2][71] + inp[72] * layer_1_weights[2][72] + inp[73] * layer_1_weights[2][73] + inp[74] * layer_1_weights[2][74] + inp[75] * layer_1_weights[2][75] + inp[76] * layer_1_weights[2][76] + inp[77] * layer_1_weights[2][77] + inp[78] * layer_1_weights[2][78] + inp[79] * layer_1_weights[2][79] + inp[80] * layer_1_weights[2][80] + inp[81] * layer_1_weights[2][81] + inp[82] * layer_1_weights[2][82] + inp[83] * layer_1_weights[2][83] + inp[84] * layer_1_weights[2][84] + inp[85] * layer_1_weights[2][85] + inp[86] * layer_1_weights[2][86] + inp[87] * layer_1_weights[2][87] + inp[88] * layer_1_weights[2][88] + inp[89] * layer_1_weights[2][89] + inp[90] * layer_1_weights[2][90] + inp[91] * layer_1_weights[2][91] + inp[92] * layer_1_weights[2][92] + inp[93] * layer_1_weights[2][93] + inp[94] * layer_1_weights[2][94] + inp[95] * layer_1_weights[2][95] + inp[96] * layer_1_weights[2][96] + inp[97] * layer_1_weights[2][97] + inp[98] * layer_1_weights[2][98] + inp[99] * layer_1_weights[2][99] + inp[100] * layer_1_weights[2][100] + inp[101] * layer_1_weights[2][101] + inp[102] * layer_1_weights[2][102] + inp[103] * layer_1_weights[2][103] + inp[104] * layer_1_weights[2][104] + inp[105] * layer_1_weights[2][105] + inp[106] * layer_1_weights[2][106] + inp[107] * layer_1_weights[2][107] + inp[108] * layer_1_weights[2][108] + inp[109] * layer_1_weights[2][109] + inp[110] * layer_1_weights[2][110] + inp[111] * layer_1_weights[2][111] + inp[112] * layer_1_weights[2][112] + inp[113] * layer_1_weights[2][113] + inp[114] * layer_1_weights[2][114] + inp[115] * layer_1_weights[2][115] + inp[116] * layer_1_weights[2][116] + inp[117] * layer_1_weights[2][117] + inp[118] * layer_1_weights[2][118] + inp[119] * layer_1_weights[2][119] + inp[120] * layer_1_weights[2][120] + inp[121] * layer_1_weights[2][121] + inp[122] * layer_1_weights[2][122] + inp[123] * layer_1_weights[2][123] + inp[124] * layer_1_weights[2][124] + inp[125] * layer_1_weights[2][125] + inp[126] * layer_1_weights[2][126] + inp[127] * layer_1_weights[2][127] + inp[128] * layer_1_weights[2][128] + inp[129] * layer_1_weights[2][129] + inp[130] * layer_1_weights[2][130] + inp[131] * layer_1_weights[2][131] + inp[132] * layer_1_weights[2][132] + inp[133] * layer_1_weights[2][133] + inp[134] * layer_1_weights[2][134] + inp[135] * layer_1_weights[2][135] + inp[136] * layer_1_weights[2][136] + inp[137] * layer_1_weights[2][137] + inp[138] * layer_1_weights[2][138] + inp[139] * layer_1_weights[2][139] + inp[140] * layer_1_weights[2][140] + inp[141] * layer_1_weights[2][141] + inp[142] * layer_1_weights[2][142] + inp[143] * layer_1_weights[2][143]);
    assign layer_1_output_3 = relu(layer_1_biases[3] + inp[0] * layer_1_weights[3][0] + inp[1] * layer_1_weights[3][1] + inp[2] * layer_1_weights[3][2] + inp[3] * layer_1_weights[3][3] + inp[4] * layer_1_weights[3][4] + inp[5] * layer_1_weights[3][5] + inp[6] * layer_1_weights[3][6] + inp[7] * layer_1_weights[3][7] + inp[8] * layer_1_weights[3][8] + inp[9] * layer_1_weights[3][9] + inp[10] * layer_1_weights[3][10] + inp[11] * layer_1_weights[3][11] + inp[12] * layer_1_weights[3][12] + inp[13] * layer_1_weights[3][13] + inp[14] * layer_1_weights[3][14] + inp[15] * layer_1_weights[3][15] + inp[16] * layer_1_weights[3][16] + inp[17] * layer_1_weights[3][17] + inp[18] * layer_1_weights[3][18] + inp[19] * layer_1_weights[3][19] + inp[20] * layer_1_weights[3][20] + inp[21] * layer_1_weights[3][21] + inp[22] * layer_1_weights[3][22] + inp[23] * layer_1_weights[3][23] + inp[24] * layer_1_weights[3][24] + inp[25] * layer_1_weights[3][25] + inp[26] * layer_1_weights[3][26] + inp[27] * layer_1_weights[3][27] + inp[28] * layer_1_weights[3][28] + inp[29] * layer_1_weights[3][29] + inp[30] * layer_1_weights[3][30] + inp[31] * layer_1_weights[3][31] + inp[32] * layer_1_weights[3][32] + inp[33] * layer_1_weights[3][33] + inp[34] * layer_1_weights[3][34] + inp[35] * layer_1_weights[3][35] + inp[36] * layer_1_weights[3][36] + inp[37] * layer_1_weights[3][37] + inp[38] * layer_1_weights[3][38] + inp[39] * layer_1_weights[3][39] + inp[40] * layer_1_weights[3][40] + inp[41] * layer_1_weights[3][41] + inp[42] * layer_1_weights[3][42] + inp[43] * layer_1_weights[3][43] + inp[44] * layer_1_weights[3][44] + inp[45] * layer_1_weights[3][45] + inp[46] * layer_1_weights[3][46] + inp[47] * layer_1_weights[3][47] + inp[48] * layer_1_weights[3][48] + inp[49] * layer_1_weights[3][49] + inp[50] * layer_1_weights[3][50] + inp[51] * layer_1_weights[3][51] + inp[52] * layer_1_weights[3][52] + inp[53] * layer_1_weights[3][53] + inp[54] * layer_1_weights[3][54] + inp[55] * layer_1_weights[3][55] + inp[56] * layer_1_weights[3][56] + inp[57] * layer_1_weights[3][57] + inp[58] * layer_1_weights[3][58] + inp[59] * layer_1_weights[3][59] + inp[60] * layer_1_weights[3][60] + inp[61] * layer_1_weights[3][61] + inp[62] * layer_1_weights[3][62] + inp[63] * layer_1_weights[3][63] + inp[64] * layer_1_weights[3][64] + inp[65] * layer_1_weights[3][65] + inp[66] * layer_1_weights[3][66] + inp[67] * layer_1_weights[3][67] + inp[68] * layer_1_weights[3][68] + inp[69] * layer_1_weights[3][69] + inp[70] * layer_1_weights[3][70] + inp[71] * layer_1_weights[3][71] + inp[72] * layer_1_weights[3][72] + inp[73] * layer_1_weights[3][73] + inp[74] * layer_1_weights[3][74] + inp[75] * layer_1_weights[3][75] + inp[76] * layer_1_weights[3][76] + inp[77] * layer_1_weights[3][77] + inp[78] * layer_1_weights[3][78] + inp[79] * layer_1_weights[3][79] + inp[80] * layer_1_weights[3][80] + inp[81] * layer_1_weights[3][81] + inp[82] * layer_1_weights[3][82] + inp[83] * layer_1_weights[3][83] + inp[84] * layer_1_weights[3][84] + inp[85] * layer_1_weights[3][85] + inp[86] * layer_1_weights[3][86] + inp[87] * layer_1_weights[3][87] + inp[88] * layer_1_weights[3][88] + inp[89] * layer_1_weights[3][89] + inp[90] * layer_1_weights[3][90] + inp[91] * layer_1_weights[3][91] + inp[92] * layer_1_weights[3][92] + inp[93] * layer_1_weights[3][93] + inp[94] * layer_1_weights[3][94] + inp[95] * layer_1_weights[3][95] + inp[96] * layer_1_weights[3][96] + inp[97] * layer_1_weights[3][97] + inp[98] * layer_1_weights[3][98] + inp[99] * layer_1_weights[3][99] + inp[100] * layer_1_weights[3][100] + inp[101] * layer_1_weights[3][101] + inp[102] * layer_1_weights[3][102] + inp[103] * layer_1_weights[3][103] + inp[104] * layer_1_weights[3][104] + inp[105] * layer_1_weights[3][105] + inp[106] * layer_1_weights[3][106] + inp[107] * layer_1_weights[3][107] + inp[108] * layer_1_weights[3][108] + inp[109] * layer_1_weights[3][109] + inp[110] * layer_1_weights[3][110] + inp[111] * layer_1_weights[3][111] + inp[112] * layer_1_weights[3][112] + inp[113] * layer_1_weights[3][113] + inp[114] * layer_1_weights[3][114] + inp[115] * layer_1_weights[3][115] + inp[116] * layer_1_weights[3][116] + inp[117] * layer_1_weights[3][117] + inp[118] * layer_1_weights[3][118] + inp[119] * layer_1_weights[3][119] + inp[120] * layer_1_weights[3][120] + inp[121] * layer_1_weights[3][121] + inp[122] * layer_1_weights[3][122] + inp[123] * layer_1_weights[3][123] + inp[124] * layer_1_weights[3][124] + inp[125] * layer_1_weights[3][125] + inp[126] * layer_1_weights[3][126] + inp[127] * layer_1_weights[3][127] + inp[128] * layer_1_weights[3][128] + inp[129] * layer_1_weights[3][129] + inp[130] * layer_1_weights[3][130] + inp[131] * layer_1_weights[3][131] + inp[132] * layer_1_weights[3][132] + inp[133] * layer_1_weights[3][133] + inp[134] * layer_1_weights[3][134] + inp[135] * layer_1_weights[3][135] + inp[136] * layer_1_weights[3][136] + inp[137] * layer_1_weights[3][137] + inp[138] * layer_1_weights[3][138] + inp[139] * layer_1_weights[3][139] + inp[140] * layer_1_weights[3][140] + inp[141] * layer_1_weights[3][141] + inp[142] * layer_1_weights[3][142] + inp[143] * layer_1_weights[3][143]);
    assign layer_1_output_4 = relu(layer_1_biases[4] + inp[0] * layer_1_weights[4][0] + inp[1] * layer_1_weights[4][1] + inp[2] * layer_1_weights[4][2] + inp[3] * layer_1_weights[4][3] + inp[4] * layer_1_weights[4][4] + inp[5] * layer_1_weights[4][5] + inp[6] * layer_1_weights[4][6] + inp[7] * layer_1_weights[4][7] + inp[8] * layer_1_weights[4][8] + inp[9] * layer_1_weights[4][9] + inp[10] * layer_1_weights[4][10] + inp[11] * layer_1_weights[4][11] + inp[12] * layer_1_weights[4][12] + inp[13] * layer_1_weights[4][13] + inp[14] * layer_1_weights[4][14] + inp[15] * layer_1_weights[4][15] + inp[16] * layer_1_weights[4][16] + inp[17] * layer_1_weights[4][17] + inp[18] * layer_1_weights[4][18] + inp[19] * layer_1_weights[4][19] + inp[20] * layer_1_weights[4][20] + inp[21] * layer_1_weights[4][21] + inp[22] * layer_1_weights[4][22] + inp[23] * layer_1_weights[4][23] + inp[24] * layer_1_weights[4][24] + inp[25] * layer_1_weights[4][25] + inp[26] * layer_1_weights[4][26] + inp[27] * layer_1_weights[4][27] + inp[28] * layer_1_weights[4][28] + inp[29] * layer_1_weights[4][29] + inp[30] * layer_1_weights[4][30] + inp[31] * layer_1_weights[4][31] + inp[32] * layer_1_weights[4][32] + inp[33] * layer_1_weights[4][33] + inp[34] * layer_1_weights[4][34] + inp[35] * layer_1_weights[4][35] + inp[36] * layer_1_weights[4][36] + inp[37] * layer_1_weights[4][37] + inp[38] * layer_1_weights[4][38] + inp[39] * layer_1_weights[4][39] + inp[40] * layer_1_weights[4][40] + inp[41] * layer_1_weights[4][41] + inp[42] * layer_1_weights[4][42] + inp[43] * layer_1_weights[4][43] + inp[44] * layer_1_weights[4][44] + inp[45] * layer_1_weights[4][45] + inp[46] * layer_1_weights[4][46] + inp[47] * layer_1_weights[4][47] + inp[48] * layer_1_weights[4][48] + inp[49] * layer_1_weights[4][49] + inp[50] * layer_1_weights[4][50] + inp[51] * layer_1_weights[4][51] + inp[52] * layer_1_weights[4][52] + inp[53] * layer_1_weights[4][53] + inp[54] * layer_1_weights[4][54] + inp[55] * layer_1_weights[4][55] + inp[56] * layer_1_weights[4][56] + inp[57] * layer_1_weights[4][57] + inp[58] * layer_1_weights[4][58] + inp[59] * layer_1_weights[4][59] + inp[60] * layer_1_weights[4][60] + inp[61] * layer_1_weights[4][61] + inp[62] * layer_1_weights[4][62] + inp[63] * layer_1_weights[4][63] + inp[64] * layer_1_weights[4][64] + inp[65] * layer_1_weights[4][65] + inp[66] * layer_1_weights[4][66] + inp[67] * layer_1_weights[4][67] + inp[68] * layer_1_weights[4][68] + inp[69] * layer_1_weights[4][69] + inp[70] * layer_1_weights[4][70] + inp[71] * layer_1_weights[4][71] + inp[72] * layer_1_weights[4][72] + inp[73] * layer_1_weights[4][73] + inp[74] * layer_1_weights[4][74] + inp[75] * layer_1_weights[4][75] + inp[76] * layer_1_weights[4][76] + inp[77] * layer_1_weights[4][77] + inp[78] * layer_1_weights[4][78] + inp[79] * layer_1_weights[4][79] + inp[80] * layer_1_weights[4][80] + inp[81] * layer_1_weights[4][81] + inp[82] * layer_1_weights[4][82] + inp[83] * layer_1_weights[4][83] + inp[84] * layer_1_weights[4][84] + inp[85] * layer_1_weights[4][85] + inp[86] * layer_1_weights[4][86] + inp[87] * layer_1_weights[4][87] + inp[88] * layer_1_weights[4][88] + inp[89] * layer_1_weights[4][89] + inp[90] * layer_1_weights[4][90] + inp[91] * layer_1_weights[4][91] + inp[92] * layer_1_weights[4][92] + inp[93] * layer_1_weights[4][93] + inp[94] * layer_1_weights[4][94] + inp[95] * layer_1_weights[4][95] + inp[96] * layer_1_weights[4][96] + inp[97] * layer_1_weights[4][97] + inp[98] * layer_1_weights[4][98] + inp[99] * layer_1_weights[4][99] + inp[100] * layer_1_weights[4][100] + inp[101] * layer_1_weights[4][101] + inp[102] * layer_1_weights[4][102] + inp[103] * layer_1_weights[4][103] + inp[104] * layer_1_weights[4][104] + inp[105] * layer_1_weights[4][105] + inp[106] * layer_1_weights[4][106] + inp[107] * layer_1_weights[4][107] + inp[108] * layer_1_weights[4][108] + inp[109] * layer_1_weights[4][109] + inp[110] * layer_1_weights[4][110] + inp[111] * layer_1_weights[4][111] + inp[112] * layer_1_weights[4][112] + inp[113] * layer_1_weights[4][113] + inp[114] * layer_1_weights[4][114] + inp[115] * layer_1_weights[4][115] + inp[116] * layer_1_weights[4][116] + inp[117] * layer_1_weights[4][117] + inp[118] * layer_1_weights[4][118] + inp[119] * layer_1_weights[4][119] + inp[120] * layer_1_weights[4][120] + inp[121] * layer_1_weights[4][121] + inp[122] * layer_1_weights[4][122] + inp[123] * layer_1_weights[4][123] + inp[124] * layer_1_weights[4][124] + inp[125] * layer_1_weights[4][125] + inp[126] * layer_1_weights[4][126] + inp[127] * layer_1_weights[4][127] + inp[128] * layer_1_weights[4][128] + inp[129] * layer_1_weights[4][129] + inp[130] * layer_1_weights[4][130] + inp[131] * layer_1_weights[4][131] + inp[132] * layer_1_weights[4][132] + inp[133] * layer_1_weights[4][133] + inp[134] * layer_1_weights[4][134] + inp[135] * layer_1_weights[4][135] + inp[136] * layer_1_weights[4][136] + inp[137] * layer_1_weights[4][137] + inp[138] * layer_1_weights[4][138] + inp[139] * layer_1_weights[4][139] + inp[140] * layer_1_weights[4][140] + inp[141] * layer_1_weights[4][141] + inp[142] * layer_1_weights[4][142] + inp[143] * layer_1_weights[4][143]);
    assign layer_1_output_5 = relu(layer_1_biases[5] + inp[0] * layer_1_weights[5][0] + inp[1] * layer_1_weights[5][1] + inp[2] * layer_1_weights[5][2] + inp[3] * layer_1_weights[5][3] + inp[4] * layer_1_weights[5][4] + inp[5] * layer_1_weights[5][5] + inp[6] * layer_1_weights[5][6] + inp[7] * layer_1_weights[5][7] + inp[8] * layer_1_weights[5][8] + inp[9] * layer_1_weights[5][9] + inp[10] * layer_1_weights[5][10] + inp[11] * layer_1_weights[5][11] + inp[12] * layer_1_weights[5][12] + inp[13] * layer_1_weights[5][13] + inp[14] * layer_1_weights[5][14] + inp[15] * layer_1_weights[5][15] + inp[16] * layer_1_weights[5][16] + inp[17] * layer_1_weights[5][17] + inp[18] * layer_1_weights[5][18] + inp[19] * layer_1_weights[5][19] + inp[20] * layer_1_weights[5][20] + inp[21] * layer_1_weights[5][21] + inp[22] * layer_1_weights[5][22] + inp[23] * layer_1_weights[5][23] + inp[24] * layer_1_weights[5][24] + inp[25] * layer_1_weights[5][25] + inp[26] * layer_1_weights[5][26] + inp[27] * layer_1_weights[5][27] + inp[28] * layer_1_weights[5][28] + inp[29] * layer_1_weights[5][29] + inp[30] * layer_1_weights[5][30] + inp[31] * layer_1_weights[5][31] + inp[32] * layer_1_weights[5][32] + inp[33] * layer_1_weights[5][33] + inp[34] * layer_1_weights[5][34] + inp[35] * layer_1_weights[5][35] + inp[36] * layer_1_weights[5][36] + inp[37] * layer_1_weights[5][37] + inp[38] * layer_1_weights[5][38] + inp[39] * layer_1_weights[5][39] + inp[40] * layer_1_weights[5][40] + inp[41] * layer_1_weights[5][41] + inp[42] * layer_1_weights[5][42] + inp[43] * layer_1_weights[5][43] + inp[44] * layer_1_weights[5][44] + inp[45] * layer_1_weights[5][45] + inp[46] * layer_1_weights[5][46] + inp[47] * layer_1_weights[5][47] + inp[48] * layer_1_weights[5][48] + inp[49] * layer_1_weights[5][49] + inp[50] * layer_1_weights[5][50] + inp[51] * layer_1_weights[5][51] + inp[52] * layer_1_weights[5][52] + inp[53] * layer_1_weights[5][53] + inp[54] * layer_1_weights[5][54] + inp[55] * layer_1_weights[5][55] + inp[56] * layer_1_weights[5][56] + inp[57] * layer_1_weights[5][57] + inp[58] * layer_1_weights[5][58] + inp[59] * layer_1_weights[5][59] + inp[60] * layer_1_weights[5][60] + inp[61] * layer_1_weights[5][61] + inp[62] * layer_1_weights[5][62] + inp[63] * layer_1_weights[5][63] + inp[64] * layer_1_weights[5][64] + inp[65] * layer_1_weights[5][65] + inp[66] * layer_1_weights[5][66] + inp[67] * layer_1_weights[5][67] + inp[68] * layer_1_weights[5][68] + inp[69] * layer_1_weights[5][69] + inp[70] * layer_1_weights[5][70] + inp[71] * layer_1_weights[5][71] + inp[72] * layer_1_weights[5][72] + inp[73] * layer_1_weights[5][73] + inp[74] * layer_1_weights[5][74] + inp[75] * layer_1_weights[5][75] + inp[76] * layer_1_weights[5][76] + inp[77] * layer_1_weights[5][77] + inp[78] * layer_1_weights[5][78] + inp[79] * layer_1_weights[5][79] + inp[80] * layer_1_weights[5][80] + inp[81] * layer_1_weights[5][81] + inp[82] * layer_1_weights[5][82] + inp[83] * layer_1_weights[5][83] + inp[84] * layer_1_weights[5][84] + inp[85] * layer_1_weights[5][85] + inp[86] * layer_1_weights[5][86] + inp[87] * layer_1_weights[5][87] + inp[88] * layer_1_weights[5][88] + inp[89] * layer_1_weights[5][89] + inp[90] * layer_1_weights[5][90] + inp[91] * layer_1_weights[5][91] + inp[92] * layer_1_weights[5][92] + inp[93] * layer_1_weights[5][93] + inp[94] * layer_1_weights[5][94] + inp[95] * layer_1_weights[5][95] + inp[96] * layer_1_weights[5][96] + inp[97] * layer_1_weights[5][97] + inp[98] * layer_1_weights[5][98] + inp[99] * layer_1_weights[5][99] + inp[100] * layer_1_weights[5][100] + inp[101] * layer_1_weights[5][101] + inp[102] * layer_1_weights[5][102] + inp[103] * layer_1_weights[5][103] + inp[104] * layer_1_weights[5][104] + inp[105] * layer_1_weights[5][105] + inp[106] * layer_1_weights[5][106] + inp[107] * layer_1_weights[5][107] + inp[108] * layer_1_weights[5][108] + inp[109] * layer_1_weights[5][109] + inp[110] * layer_1_weights[5][110] + inp[111] * layer_1_weights[5][111] + inp[112] * layer_1_weights[5][112] + inp[113] * layer_1_weights[5][113] + inp[114] * layer_1_weights[5][114] + inp[115] * layer_1_weights[5][115] + inp[116] * layer_1_weights[5][116] + inp[117] * layer_1_weights[5][117] + inp[118] * layer_1_weights[5][118] + inp[119] * layer_1_weights[5][119] + inp[120] * layer_1_weights[5][120] + inp[121] * layer_1_weights[5][121] + inp[122] * layer_1_weights[5][122] + inp[123] * layer_1_weights[5][123] + inp[124] * layer_1_weights[5][124] + inp[125] * layer_1_weights[5][125] + inp[126] * layer_1_weights[5][126] + inp[127] * layer_1_weights[5][127] + inp[128] * layer_1_weights[5][128] + inp[129] * layer_1_weights[5][129] + inp[130] * layer_1_weights[5][130] + inp[131] * layer_1_weights[5][131] + inp[132] * layer_1_weights[5][132] + inp[133] * layer_1_weights[5][133] + inp[134] * layer_1_weights[5][134] + inp[135] * layer_1_weights[5][135] + inp[136] * layer_1_weights[5][136] + inp[137] * layer_1_weights[5][137] + inp[138] * layer_1_weights[5][138] + inp[139] * layer_1_weights[5][139] + inp[140] * layer_1_weights[5][140] + inp[141] * layer_1_weights[5][141] + inp[142] * layer_1_weights[5][142] + inp[143] * layer_1_weights[5][143]);
    assign layer_1_output_6 = relu(layer_1_biases[6] + inp[0] * layer_1_weights[6][0] + inp[1] * layer_1_weights[6][1] + inp[2] * layer_1_weights[6][2] + inp[3] * layer_1_weights[6][3] + inp[4] * layer_1_weights[6][4] + inp[5] * layer_1_weights[6][5] + inp[6] * layer_1_weights[6][6] + inp[7] * layer_1_weights[6][7] + inp[8] * layer_1_weights[6][8] + inp[9] * layer_1_weights[6][9] + inp[10] * layer_1_weights[6][10] + inp[11] * layer_1_weights[6][11] + inp[12] * layer_1_weights[6][12] + inp[13] * layer_1_weights[6][13] + inp[14] * layer_1_weights[6][14] + inp[15] * layer_1_weights[6][15] + inp[16] * layer_1_weights[6][16] + inp[17] * layer_1_weights[6][17] + inp[18] * layer_1_weights[6][18] + inp[19] * layer_1_weights[6][19] + inp[20] * layer_1_weights[6][20] + inp[21] * layer_1_weights[6][21] + inp[22] * layer_1_weights[6][22] + inp[23] * layer_1_weights[6][23] + inp[24] * layer_1_weights[6][24] + inp[25] * layer_1_weights[6][25] + inp[26] * layer_1_weights[6][26] + inp[27] * layer_1_weights[6][27] + inp[28] * layer_1_weights[6][28] + inp[29] * layer_1_weights[6][29] + inp[30] * layer_1_weights[6][30] + inp[31] * layer_1_weights[6][31] + inp[32] * layer_1_weights[6][32] + inp[33] * layer_1_weights[6][33] + inp[34] * layer_1_weights[6][34] + inp[35] * layer_1_weights[6][35] + inp[36] * layer_1_weights[6][36] + inp[37] * layer_1_weights[6][37] + inp[38] * layer_1_weights[6][38] + inp[39] * layer_1_weights[6][39] + inp[40] * layer_1_weights[6][40] + inp[41] * layer_1_weights[6][41] + inp[42] * layer_1_weights[6][42] + inp[43] * layer_1_weights[6][43] + inp[44] * layer_1_weights[6][44] + inp[45] * layer_1_weights[6][45] + inp[46] * layer_1_weights[6][46] + inp[47] * layer_1_weights[6][47] + inp[48] * layer_1_weights[6][48] + inp[49] * layer_1_weights[6][49] + inp[50] * layer_1_weights[6][50] + inp[51] * layer_1_weights[6][51] + inp[52] * layer_1_weights[6][52] + inp[53] * layer_1_weights[6][53] + inp[54] * layer_1_weights[6][54] + inp[55] * layer_1_weights[6][55] + inp[56] * layer_1_weights[6][56] + inp[57] * layer_1_weights[6][57] + inp[58] * layer_1_weights[6][58] + inp[59] * layer_1_weights[6][59] + inp[60] * layer_1_weights[6][60] + inp[61] * layer_1_weights[6][61] + inp[62] * layer_1_weights[6][62] + inp[63] * layer_1_weights[6][63] + inp[64] * layer_1_weights[6][64] + inp[65] * layer_1_weights[6][65] + inp[66] * layer_1_weights[6][66] + inp[67] * layer_1_weights[6][67] + inp[68] * layer_1_weights[6][68] + inp[69] * layer_1_weights[6][69] + inp[70] * layer_1_weights[6][70] + inp[71] * layer_1_weights[6][71] + inp[72] * layer_1_weights[6][72] + inp[73] * layer_1_weights[6][73] + inp[74] * layer_1_weights[6][74] + inp[75] * layer_1_weights[6][75] + inp[76] * layer_1_weights[6][76] + inp[77] * layer_1_weights[6][77] + inp[78] * layer_1_weights[6][78] + inp[79] * layer_1_weights[6][79] + inp[80] * layer_1_weights[6][80] + inp[81] * layer_1_weights[6][81] + inp[82] * layer_1_weights[6][82] + inp[83] * layer_1_weights[6][83] + inp[84] * layer_1_weights[6][84] + inp[85] * layer_1_weights[6][85] + inp[86] * layer_1_weights[6][86] + inp[87] * layer_1_weights[6][87] + inp[88] * layer_1_weights[6][88] + inp[89] * layer_1_weights[6][89] + inp[90] * layer_1_weights[6][90] + inp[91] * layer_1_weights[6][91] + inp[92] * layer_1_weights[6][92] + inp[93] * layer_1_weights[6][93] + inp[94] * layer_1_weights[6][94] + inp[95] * layer_1_weights[6][95] + inp[96] * layer_1_weights[6][96] + inp[97] * layer_1_weights[6][97] + inp[98] * layer_1_weights[6][98] + inp[99] * layer_1_weights[6][99] + inp[100] * layer_1_weights[6][100] + inp[101] * layer_1_weights[6][101] + inp[102] * layer_1_weights[6][102] + inp[103] * layer_1_weights[6][103] + inp[104] * layer_1_weights[6][104] + inp[105] * layer_1_weights[6][105] + inp[106] * layer_1_weights[6][106] + inp[107] * layer_1_weights[6][107] + inp[108] * layer_1_weights[6][108] + inp[109] * layer_1_weights[6][109] + inp[110] * layer_1_weights[6][110] + inp[111] * layer_1_weights[6][111] + inp[112] * layer_1_weights[6][112] + inp[113] * layer_1_weights[6][113] + inp[114] * layer_1_weights[6][114] + inp[115] * layer_1_weights[6][115] + inp[116] * layer_1_weights[6][116] + inp[117] * layer_1_weights[6][117] + inp[118] * layer_1_weights[6][118] + inp[119] * layer_1_weights[6][119] + inp[120] * layer_1_weights[6][120] + inp[121] * layer_1_weights[6][121] + inp[122] * layer_1_weights[6][122] + inp[123] * layer_1_weights[6][123] + inp[124] * layer_1_weights[6][124] + inp[125] * layer_1_weights[6][125] + inp[126] * layer_1_weights[6][126] + inp[127] * layer_1_weights[6][127] + inp[128] * layer_1_weights[6][128] + inp[129] * layer_1_weights[6][129] + inp[130] * layer_1_weights[6][130] + inp[131] * layer_1_weights[6][131] + inp[132] * layer_1_weights[6][132] + inp[133] * layer_1_weights[6][133] + inp[134] * layer_1_weights[6][134] + inp[135] * layer_1_weights[6][135] + inp[136] * layer_1_weights[6][136] + inp[137] * layer_1_weights[6][137] + inp[138] * layer_1_weights[6][138] + inp[139] * layer_1_weights[6][139] + inp[140] * layer_1_weights[6][140] + inp[141] * layer_1_weights[6][141] + inp[142] * layer_1_weights[6][142] + inp[143] * layer_1_weights[6][143]);
    assign layer_1_output_7 = relu(layer_1_biases[7] + inp[0] * layer_1_weights[7][0] + inp[1] * layer_1_weights[7][1] + inp[2] * layer_1_weights[7][2] + inp[3] * layer_1_weights[7][3] + inp[4] * layer_1_weights[7][4] + inp[5] * layer_1_weights[7][5] + inp[6] * layer_1_weights[7][6] + inp[7] * layer_1_weights[7][7] + inp[8] * layer_1_weights[7][8] + inp[9] * layer_1_weights[7][9] + inp[10] * layer_1_weights[7][10] + inp[11] * layer_1_weights[7][11] + inp[12] * layer_1_weights[7][12] + inp[13] * layer_1_weights[7][13] + inp[14] * layer_1_weights[7][14] + inp[15] * layer_1_weights[7][15] + inp[16] * layer_1_weights[7][16] + inp[17] * layer_1_weights[7][17] + inp[18] * layer_1_weights[7][18] + inp[19] * layer_1_weights[7][19] + inp[20] * layer_1_weights[7][20] + inp[21] * layer_1_weights[7][21] + inp[22] * layer_1_weights[7][22] + inp[23] * layer_1_weights[7][23] + inp[24] * layer_1_weights[7][24] + inp[25] * layer_1_weights[7][25] + inp[26] * layer_1_weights[7][26] + inp[27] * layer_1_weights[7][27] + inp[28] * layer_1_weights[7][28] + inp[29] * layer_1_weights[7][29] + inp[30] * layer_1_weights[7][30] + inp[31] * layer_1_weights[7][31] + inp[32] * layer_1_weights[7][32] + inp[33] * layer_1_weights[7][33] + inp[34] * layer_1_weights[7][34] + inp[35] * layer_1_weights[7][35] + inp[36] * layer_1_weights[7][36] + inp[37] * layer_1_weights[7][37] + inp[38] * layer_1_weights[7][38] + inp[39] * layer_1_weights[7][39] + inp[40] * layer_1_weights[7][40] + inp[41] * layer_1_weights[7][41] + inp[42] * layer_1_weights[7][42] + inp[43] * layer_1_weights[7][43] + inp[44] * layer_1_weights[7][44] + inp[45] * layer_1_weights[7][45] + inp[46] * layer_1_weights[7][46] + inp[47] * layer_1_weights[7][47] + inp[48] * layer_1_weights[7][48] + inp[49] * layer_1_weights[7][49] + inp[50] * layer_1_weights[7][50] + inp[51] * layer_1_weights[7][51] + inp[52] * layer_1_weights[7][52] + inp[53] * layer_1_weights[7][53] + inp[54] * layer_1_weights[7][54] + inp[55] * layer_1_weights[7][55] + inp[56] * layer_1_weights[7][56] + inp[57] * layer_1_weights[7][57] + inp[58] * layer_1_weights[7][58] + inp[59] * layer_1_weights[7][59] + inp[60] * layer_1_weights[7][60] + inp[61] * layer_1_weights[7][61] + inp[62] * layer_1_weights[7][62] + inp[63] * layer_1_weights[7][63] + inp[64] * layer_1_weights[7][64] + inp[65] * layer_1_weights[7][65] + inp[66] * layer_1_weights[7][66] + inp[67] * layer_1_weights[7][67] + inp[68] * layer_1_weights[7][68] + inp[69] * layer_1_weights[7][69] + inp[70] * layer_1_weights[7][70] + inp[71] * layer_1_weights[7][71] + inp[72] * layer_1_weights[7][72] + inp[73] * layer_1_weights[7][73] + inp[74] * layer_1_weights[7][74] + inp[75] * layer_1_weights[7][75] + inp[76] * layer_1_weights[7][76] + inp[77] * layer_1_weights[7][77] + inp[78] * layer_1_weights[7][78] + inp[79] * layer_1_weights[7][79] + inp[80] * layer_1_weights[7][80] + inp[81] * layer_1_weights[7][81] + inp[82] * layer_1_weights[7][82] + inp[83] * layer_1_weights[7][83] + inp[84] * layer_1_weights[7][84] + inp[85] * layer_1_weights[7][85] + inp[86] * layer_1_weights[7][86] + inp[87] * layer_1_weights[7][87] + inp[88] * layer_1_weights[7][88] + inp[89] * layer_1_weights[7][89] + inp[90] * layer_1_weights[7][90] + inp[91] * layer_1_weights[7][91] + inp[92] * layer_1_weights[7][92] + inp[93] * layer_1_weights[7][93] + inp[94] * layer_1_weights[7][94] + inp[95] * layer_1_weights[7][95] + inp[96] * layer_1_weights[7][96] + inp[97] * layer_1_weights[7][97] + inp[98] * layer_1_weights[7][98] + inp[99] * layer_1_weights[7][99] + inp[100] * layer_1_weights[7][100] + inp[101] * layer_1_weights[7][101] + inp[102] * layer_1_weights[7][102] + inp[103] * layer_1_weights[7][103] + inp[104] * layer_1_weights[7][104] + inp[105] * layer_1_weights[7][105] + inp[106] * layer_1_weights[7][106] + inp[107] * layer_1_weights[7][107] + inp[108] * layer_1_weights[7][108] + inp[109] * layer_1_weights[7][109] + inp[110] * layer_1_weights[7][110] + inp[111] * layer_1_weights[7][111] + inp[112] * layer_1_weights[7][112] + inp[113] * layer_1_weights[7][113] + inp[114] * layer_1_weights[7][114] + inp[115] * layer_1_weights[7][115] + inp[116] * layer_1_weights[7][116] + inp[117] * layer_1_weights[7][117] + inp[118] * layer_1_weights[7][118] + inp[119] * layer_1_weights[7][119] + inp[120] * layer_1_weights[7][120] + inp[121] * layer_1_weights[7][121] + inp[122] * layer_1_weights[7][122] + inp[123] * layer_1_weights[7][123] + inp[124] * layer_1_weights[7][124] + inp[125] * layer_1_weights[7][125] + inp[126] * layer_1_weights[7][126] + inp[127] * layer_1_weights[7][127] + inp[128] * layer_1_weights[7][128] + inp[129] * layer_1_weights[7][129] + inp[130] * layer_1_weights[7][130] + inp[131] * layer_1_weights[7][131] + inp[132] * layer_1_weights[7][132] + inp[133] * layer_1_weights[7][133] + inp[134] * layer_1_weights[7][134] + inp[135] * layer_1_weights[7][135] + inp[136] * layer_1_weights[7][136] + inp[137] * layer_1_weights[7][137] + inp[138] * layer_1_weights[7][138] + inp[139] * layer_1_weights[7][139] + inp[140] * layer_1_weights[7][140] + inp[141] * layer_1_weights[7][141] + inp[142] * layer_1_weights[7][142] + inp[143] * layer_1_weights[7][143]);
    assign layer_1_output_8 = relu(layer_1_biases[8] + inp[0] * layer_1_weights[8][0] + inp[1] * layer_1_weights[8][1] + inp[2] * layer_1_weights[8][2] + inp[3] * layer_1_weights[8][3] + inp[4] * layer_1_weights[8][4] + inp[5] * layer_1_weights[8][5] + inp[6] * layer_1_weights[8][6] + inp[7] * layer_1_weights[8][7] + inp[8] * layer_1_weights[8][8] + inp[9] * layer_1_weights[8][9] + inp[10] * layer_1_weights[8][10] + inp[11] * layer_1_weights[8][11] + inp[12] * layer_1_weights[8][12] + inp[13] * layer_1_weights[8][13] + inp[14] * layer_1_weights[8][14] + inp[15] * layer_1_weights[8][15] + inp[16] * layer_1_weights[8][16] + inp[17] * layer_1_weights[8][17] + inp[18] * layer_1_weights[8][18] + inp[19] * layer_1_weights[8][19] + inp[20] * layer_1_weights[8][20] + inp[21] * layer_1_weights[8][21] + inp[22] * layer_1_weights[8][22] + inp[23] * layer_1_weights[8][23] + inp[24] * layer_1_weights[8][24] + inp[25] * layer_1_weights[8][25] + inp[26] * layer_1_weights[8][26] + inp[27] * layer_1_weights[8][27] + inp[28] * layer_1_weights[8][28] + inp[29] * layer_1_weights[8][29] + inp[30] * layer_1_weights[8][30] + inp[31] * layer_1_weights[8][31] + inp[32] * layer_1_weights[8][32] + inp[33] * layer_1_weights[8][33] + inp[34] * layer_1_weights[8][34] + inp[35] * layer_1_weights[8][35] + inp[36] * layer_1_weights[8][36] + inp[37] * layer_1_weights[8][37] + inp[38] * layer_1_weights[8][38] + inp[39] * layer_1_weights[8][39] + inp[40] * layer_1_weights[8][40] + inp[41] * layer_1_weights[8][41] + inp[42] * layer_1_weights[8][42] + inp[43] * layer_1_weights[8][43] + inp[44] * layer_1_weights[8][44] + inp[45] * layer_1_weights[8][45] + inp[46] * layer_1_weights[8][46] + inp[47] * layer_1_weights[8][47] + inp[48] * layer_1_weights[8][48] + inp[49] * layer_1_weights[8][49] + inp[50] * layer_1_weights[8][50] + inp[51] * layer_1_weights[8][51] + inp[52] * layer_1_weights[8][52] + inp[53] * layer_1_weights[8][53] + inp[54] * layer_1_weights[8][54] + inp[55] * layer_1_weights[8][55] + inp[56] * layer_1_weights[8][56] + inp[57] * layer_1_weights[8][57] + inp[58] * layer_1_weights[8][58] + inp[59] * layer_1_weights[8][59] + inp[60] * layer_1_weights[8][60] + inp[61] * layer_1_weights[8][61] + inp[62] * layer_1_weights[8][62] + inp[63] * layer_1_weights[8][63] + inp[64] * layer_1_weights[8][64] + inp[65] * layer_1_weights[8][65] + inp[66] * layer_1_weights[8][66] + inp[67] * layer_1_weights[8][67] + inp[68] * layer_1_weights[8][68] + inp[69] * layer_1_weights[8][69] + inp[70] * layer_1_weights[8][70] + inp[71] * layer_1_weights[8][71] + inp[72] * layer_1_weights[8][72] + inp[73] * layer_1_weights[8][73] + inp[74] * layer_1_weights[8][74] + inp[75] * layer_1_weights[8][75] + inp[76] * layer_1_weights[8][76] + inp[77] * layer_1_weights[8][77] + inp[78] * layer_1_weights[8][78] + inp[79] * layer_1_weights[8][79] + inp[80] * layer_1_weights[8][80] + inp[81] * layer_1_weights[8][81] + inp[82] * layer_1_weights[8][82] + inp[83] * layer_1_weights[8][83] + inp[84] * layer_1_weights[8][84] + inp[85] * layer_1_weights[8][85] + inp[86] * layer_1_weights[8][86] + inp[87] * layer_1_weights[8][87] + inp[88] * layer_1_weights[8][88] + inp[89] * layer_1_weights[8][89] + inp[90] * layer_1_weights[8][90] + inp[91] * layer_1_weights[8][91] + inp[92] * layer_1_weights[8][92] + inp[93] * layer_1_weights[8][93] + inp[94] * layer_1_weights[8][94] + inp[95] * layer_1_weights[8][95] + inp[96] * layer_1_weights[8][96] + inp[97] * layer_1_weights[8][97] + inp[98] * layer_1_weights[8][98] + inp[99] * layer_1_weights[8][99] + inp[100] * layer_1_weights[8][100] + inp[101] * layer_1_weights[8][101] + inp[102] * layer_1_weights[8][102] + inp[103] * layer_1_weights[8][103] + inp[104] * layer_1_weights[8][104] + inp[105] * layer_1_weights[8][105] + inp[106] * layer_1_weights[8][106] + inp[107] * layer_1_weights[8][107] + inp[108] * layer_1_weights[8][108] + inp[109] * layer_1_weights[8][109] + inp[110] * layer_1_weights[8][110] + inp[111] * layer_1_weights[8][111] + inp[112] * layer_1_weights[8][112] + inp[113] * layer_1_weights[8][113] + inp[114] * layer_1_weights[8][114] + inp[115] * layer_1_weights[8][115] + inp[116] * layer_1_weights[8][116] + inp[117] * layer_1_weights[8][117] + inp[118] * layer_1_weights[8][118] + inp[119] * layer_1_weights[8][119] + inp[120] * layer_1_weights[8][120] + inp[121] * layer_1_weights[8][121] + inp[122] * layer_1_weights[8][122] + inp[123] * layer_1_weights[8][123] + inp[124] * layer_1_weights[8][124] + inp[125] * layer_1_weights[8][125] + inp[126] * layer_1_weights[8][126] + inp[127] * layer_1_weights[8][127] + inp[128] * layer_1_weights[8][128] + inp[129] * layer_1_weights[8][129] + inp[130] * layer_1_weights[8][130] + inp[131] * layer_1_weights[8][131] + inp[132] * layer_1_weights[8][132] + inp[133] * layer_1_weights[8][133] + inp[134] * layer_1_weights[8][134] + inp[135] * layer_1_weights[8][135] + inp[136] * layer_1_weights[8][136] + inp[137] * layer_1_weights[8][137] + inp[138] * layer_1_weights[8][138] + inp[139] * layer_1_weights[8][139] + inp[140] * layer_1_weights[8][140] + inp[141] * layer_1_weights[8][141] + inp[142] * layer_1_weights[8][142] + inp[143] * layer_1_weights[8][143]);
    assign layer_1_output_9 = relu(layer_1_biases[9] + inp[0] * layer_1_weights[9][0] + inp[1] * layer_1_weights[9][1] + inp[2] * layer_1_weights[9][2] + inp[3] * layer_1_weights[9][3] + inp[4] * layer_1_weights[9][4] + inp[5] * layer_1_weights[9][5] + inp[6] * layer_1_weights[9][6] + inp[7] * layer_1_weights[9][7] + inp[8] * layer_1_weights[9][8] + inp[9] * layer_1_weights[9][9] + inp[10] * layer_1_weights[9][10] + inp[11] * layer_1_weights[9][11] + inp[12] * layer_1_weights[9][12] + inp[13] * layer_1_weights[9][13] + inp[14] * layer_1_weights[9][14] + inp[15] * layer_1_weights[9][15] + inp[16] * layer_1_weights[9][16] + inp[17] * layer_1_weights[9][17] + inp[18] * layer_1_weights[9][18] + inp[19] * layer_1_weights[9][19] + inp[20] * layer_1_weights[9][20] + inp[21] * layer_1_weights[9][21] + inp[22] * layer_1_weights[9][22] + inp[23] * layer_1_weights[9][23] + inp[24] * layer_1_weights[9][24] + inp[25] * layer_1_weights[9][25] + inp[26] * layer_1_weights[9][26] + inp[27] * layer_1_weights[9][27] + inp[28] * layer_1_weights[9][28] + inp[29] * layer_1_weights[9][29] + inp[30] * layer_1_weights[9][30] + inp[31] * layer_1_weights[9][31] + inp[32] * layer_1_weights[9][32] + inp[33] * layer_1_weights[9][33] + inp[34] * layer_1_weights[9][34] + inp[35] * layer_1_weights[9][35] + inp[36] * layer_1_weights[9][36] + inp[37] * layer_1_weights[9][37] + inp[38] * layer_1_weights[9][38] + inp[39] * layer_1_weights[9][39] + inp[40] * layer_1_weights[9][40] + inp[41] * layer_1_weights[9][41] + inp[42] * layer_1_weights[9][42] + inp[43] * layer_1_weights[9][43] + inp[44] * layer_1_weights[9][44] + inp[45] * layer_1_weights[9][45] + inp[46] * layer_1_weights[9][46] + inp[47] * layer_1_weights[9][47] + inp[48] * layer_1_weights[9][48] + inp[49] * layer_1_weights[9][49] + inp[50] * layer_1_weights[9][50] + inp[51] * layer_1_weights[9][51] + inp[52] * layer_1_weights[9][52] + inp[53] * layer_1_weights[9][53] + inp[54] * layer_1_weights[9][54] + inp[55] * layer_1_weights[9][55] + inp[56] * layer_1_weights[9][56] + inp[57] * layer_1_weights[9][57] + inp[58] * layer_1_weights[9][58] + inp[59] * layer_1_weights[9][59] + inp[60] * layer_1_weights[9][60] + inp[61] * layer_1_weights[9][61] + inp[62] * layer_1_weights[9][62] + inp[63] * layer_1_weights[9][63] + inp[64] * layer_1_weights[9][64] + inp[65] * layer_1_weights[9][65] + inp[66] * layer_1_weights[9][66] + inp[67] * layer_1_weights[9][67] + inp[68] * layer_1_weights[9][68] + inp[69] * layer_1_weights[9][69] + inp[70] * layer_1_weights[9][70] + inp[71] * layer_1_weights[9][71] + inp[72] * layer_1_weights[9][72] + inp[73] * layer_1_weights[9][73] + inp[74] * layer_1_weights[9][74] + inp[75] * layer_1_weights[9][75] + inp[76] * layer_1_weights[9][76] + inp[77] * layer_1_weights[9][77] + inp[78] * layer_1_weights[9][78] + inp[79] * layer_1_weights[9][79] + inp[80] * layer_1_weights[9][80] + inp[81] * layer_1_weights[9][81] + inp[82] * layer_1_weights[9][82] + inp[83] * layer_1_weights[9][83] + inp[84] * layer_1_weights[9][84] + inp[85] * layer_1_weights[9][85] + inp[86] * layer_1_weights[9][86] + inp[87] * layer_1_weights[9][87] + inp[88] * layer_1_weights[9][88] + inp[89] * layer_1_weights[9][89] + inp[90] * layer_1_weights[9][90] + inp[91] * layer_1_weights[9][91] + inp[92] * layer_1_weights[9][92] + inp[93] * layer_1_weights[9][93] + inp[94] * layer_1_weights[9][94] + inp[95] * layer_1_weights[9][95] + inp[96] * layer_1_weights[9][96] + inp[97] * layer_1_weights[9][97] + inp[98] * layer_1_weights[9][98] + inp[99] * layer_1_weights[9][99] + inp[100] * layer_1_weights[9][100] + inp[101] * layer_1_weights[9][101] + inp[102] * layer_1_weights[9][102] + inp[103] * layer_1_weights[9][103] + inp[104] * layer_1_weights[9][104] + inp[105] * layer_1_weights[9][105] + inp[106] * layer_1_weights[9][106] + inp[107] * layer_1_weights[9][107] + inp[108] * layer_1_weights[9][108] + inp[109] * layer_1_weights[9][109] + inp[110] * layer_1_weights[9][110] + inp[111] * layer_1_weights[9][111] + inp[112] * layer_1_weights[9][112] + inp[113] * layer_1_weights[9][113] + inp[114] * layer_1_weights[9][114] + inp[115] * layer_1_weights[9][115] + inp[116] * layer_1_weights[9][116] + inp[117] * layer_1_weights[9][117] + inp[118] * layer_1_weights[9][118] + inp[119] * layer_1_weights[9][119] + inp[120] * layer_1_weights[9][120] + inp[121] * layer_1_weights[9][121] + inp[122] * layer_1_weights[9][122] + inp[123] * layer_1_weights[9][123] + inp[124] * layer_1_weights[9][124] + inp[125] * layer_1_weights[9][125] + inp[126] * layer_1_weights[9][126] + inp[127] * layer_1_weights[9][127] + inp[128] * layer_1_weights[9][128] + inp[129] * layer_1_weights[9][129] + inp[130] * layer_1_weights[9][130] + inp[131] * layer_1_weights[9][131] + inp[132] * layer_1_weights[9][132] + inp[133] * layer_1_weights[9][133] + inp[134] * layer_1_weights[9][134] + inp[135] * layer_1_weights[9][135] + inp[136] * layer_1_weights[9][136] + inp[137] * layer_1_weights[9][137] + inp[138] * layer_1_weights[9][138] + inp[139] * layer_1_weights[9][139] + inp[140] * layer_1_weights[9][140] + inp[141] * layer_1_weights[9][141] + inp[142] * layer_1_weights[9][142] + inp[143] * layer_1_weights[9][143]);
    assign layer_1_output_10 = relu(layer_1_biases[10] + inp[0] * layer_1_weights[10][0] + inp[1] * layer_1_weights[10][1] + inp[2] * layer_1_weights[10][2] + inp[3] * layer_1_weights[10][3] + inp[4] * layer_1_weights[10][4] + inp[5] * layer_1_weights[10][5] + inp[6] * layer_1_weights[10][6] + inp[7] * layer_1_weights[10][7] + inp[8] * layer_1_weights[10][8] + inp[9] * layer_1_weights[10][9] + inp[10] * layer_1_weights[10][10] + inp[11] * layer_1_weights[10][11] + inp[12] * layer_1_weights[10][12] + inp[13] * layer_1_weights[10][13] + inp[14] * layer_1_weights[10][14] + inp[15] * layer_1_weights[10][15] + inp[16] * layer_1_weights[10][16] + inp[17] * layer_1_weights[10][17] + inp[18] * layer_1_weights[10][18] + inp[19] * layer_1_weights[10][19] + inp[20] * layer_1_weights[10][20] + inp[21] * layer_1_weights[10][21] + inp[22] * layer_1_weights[10][22] + inp[23] * layer_1_weights[10][23] + inp[24] * layer_1_weights[10][24] + inp[25] * layer_1_weights[10][25] + inp[26] * layer_1_weights[10][26] + inp[27] * layer_1_weights[10][27] + inp[28] * layer_1_weights[10][28] + inp[29] * layer_1_weights[10][29] + inp[30] * layer_1_weights[10][30] + inp[31] * layer_1_weights[10][31] + inp[32] * layer_1_weights[10][32] + inp[33] * layer_1_weights[10][33] + inp[34] * layer_1_weights[10][34] + inp[35] * layer_1_weights[10][35] + inp[36] * layer_1_weights[10][36] + inp[37] * layer_1_weights[10][37] + inp[38] * layer_1_weights[10][38] + inp[39] * layer_1_weights[10][39] + inp[40] * layer_1_weights[10][40] + inp[41] * layer_1_weights[10][41] + inp[42] * layer_1_weights[10][42] + inp[43] * layer_1_weights[10][43] + inp[44] * layer_1_weights[10][44] + inp[45] * layer_1_weights[10][45] + inp[46] * layer_1_weights[10][46] + inp[47] * layer_1_weights[10][47] + inp[48] * layer_1_weights[10][48] + inp[49] * layer_1_weights[10][49] + inp[50] * layer_1_weights[10][50] + inp[51] * layer_1_weights[10][51] + inp[52] * layer_1_weights[10][52] + inp[53] * layer_1_weights[10][53] + inp[54] * layer_1_weights[10][54] + inp[55] * layer_1_weights[10][55] + inp[56] * layer_1_weights[10][56] + inp[57] * layer_1_weights[10][57] + inp[58] * layer_1_weights[10][58] + inp[59] * layer_1_weights[10][59] + inp[60] * layer_1_weights[10][60] + inp[61] * layer_1_weights[10][61] + inp[62] * layer_1_weights[10][62] + inp[63] * layer_1_weights[10][63] + inp[64] * layer_1_weights[10][64] + inp[65] * layer_1_weights[10][65] + inp[66] * layer_1_weights[10][66] + inp[67] * layer_1_weights[10][67] + inp[68] * layer_1_weights[10][68] + inp[69] * layer_1_weights[10][69] + inp[70] * layer_1_weights[10][70] + inp[71] * layer_1_weights[10][71] + inp[72] * layer_1_weights[10][72] + inp[73] * layer_1_weights[10][73] + inp[74] * layer_1_weights[10][74] + inp[75] * layer_1_weights[10][75] + inp[76] * layer_1_weights[10][76] + inp[77] * layer_1_weights[10][77] + inp[78] * layer_1_weights[10][78] + inp[79] * layer_1_weights[10][79] + inp[80] * layer_1_weights[10][80] + inp[81] * layer_1_weights[10][81] + inp[82] * layer_1_weights[10][82] + inp[83] * layer_1_weights[10][83] + inp[84] * layer_1_weights[10][84] + inp[85] * layer_1_weights[10][85] + inp[86] * layer_1_weights[10][86] + inp[87] * layer_1_weights[10][87] + inp[88] * layer_1_weights[10][88] + inp[89] * layer_1_weights[10][89] + inp[90] * layer_1_weights[10][90] + inp[91] * layer_1_weights[10][91] + inp[92] * layer_1_weights[10][92] + inp[93] * layer_1_weights[10][93] + inp[94] * layer_1_weights[10][94] + inp[95] * layer_1_weights[10][95] + inp[96] * layer_1_weights[10][96] + inp[97] * layer_1_weights[10][97] + inp[98] * layer_1_weights[10][98] + inp[99] * layer_1_weights[10][99] + inp[100] * layer_1_weights[10][100] + inp[101] * layer_1_weights[10][101] + inp[102] * layer_1_weights[10][102] + inp[103] * layer_1_weights[10][103] + inp[104] * layer_1_weights[10][104] + inp[105] * layer_1_weights[10][105] + inp[106] * layer_1_weights[10][106] + inp[107] * layer_1_weights[10][107] + inp[108] * layer_1_weights[10][108] + inp[109] * layer_1_weights[10][109] + inp[110] * layer_1_weights[10][110] + inp[111] * layer_1_weights[10][111] + inp[112] * layer_1_weights[10][112] + inp[113] * layer_1_weights[10][113] + inp[114] * layer_1_weights[10][114] + inp[115] * layer_1_weights[10][115] + inp[116] * layer_1_weights[10][116] + inp[117] * layer_1_weights[10][117] + inp[118] * layer_1_weights[10][118] + inp[119] * layer_1_weights[10][119] + inp[120] * layer_1_weights[10][120] + inp[121] * layer_1_weights[10][121] + inp[122] * layer_1_weights[10][122] + inp[123] * layer_1_weights[10][123] + inp[124] * layer_1_weights[10][124] + inp[125] * layer_1_weights[10][125] + inp[126] * layer_1_weights[10][126] + inp[127] * layer_1_weights[10][127] + inp[128] * layer_1_weights[10][128] + inp[129] * layer_1_weights[10][129] + inp[130] * layer_1_weights[10][130] + inp[131] * layer_1_weights[10][131] + inp[132] * layer_1_weights[10][132] + inp[133] * layer_1_weights[10][133] + inp[134] * layer_1_weights[10][134] + inp[135] * layer_1_weights[10][135] + inp[136] * layer_1_weights[10][136] + inp[137] * layer_1_weights[10][137] + inp[138] * layer_1_weights[10][138] + inp[139] * layer_1_weights[10][139] + inp[140] * layer_1_weights[10][140] + inp[141] * layer_1_weights[10][141] + inp[142] * layer_1_weights[10][142] + inp[143] * layer_1_weights[10][143]);
    assign layer_1_output_11 = relu(layer_1_biases[11] + inp[0] * layer_1_weights[11][0] + inp[1] * layer_1_weights[11][1] + inp[2] * layer_1_weights[11][2] + inp[3] * layer_1_weights[11][3] + inp[4] * layer_1_weights[11][4] + inp[5] * layer_1_weights[11][5] + inp[6] * layer_1_weights[11][6] + inp[7] * layer_1_weights[11][7] + inp[8] * layer_1_weights[11][8] + inp[9] * layer_1_weights[11][9] + inp[10] * layer_1_weights[11][10] + inp[11] * layer_1_weights[11][11] + inp[12] * layer_1_weights[11][12] + inp[13] * layer_1_weights[11][13] + inp[14] * layer_1_weights[11][14] + inp[15] * layer_1_weights[11][15] + inp[16] * layer_1_weights[11][16] + inp[17] * layer_1_weights[11][17] + inp[18] * layer_1_weights[11][18] + inp[19] * layer_1_weights[11][19] + inp[20] * layer_1_weights[11][20] + inp[21] * layer_1_weights[11][21] + inp[22] * layer_1_weights[11][22] + inp[23] * layer_1_weights[11][23] + inp[24] * layer_1_weights[11][24] + inp[25] * layer_1_weights[11][25] + inp[26] * layer_1_weights[11][26] + inp[27] * layer_1_weights[11][27] + inp[28] * layer_1_weights[11][28] + inp[29] * layer_1_weights[11][29] + inp[30] * layer_1_weights[11][30] + inp[31] * layer_1_weights[11][31] + inp[32] * layer_1_weights[11][32] + inp[33] * layer_1_weights[11][33] + inp[34] * layer_1_weights[11][34] + inp[35] * layer_1_weights[11][35] + inp[36] * layer_1_weights[11][36] + inp[37] * layer_1_weights[11][37] + inp[38] * layer_1_weights[11][38] + inp[39] * layer_1_weights[11][39] + inp[40] * layer_1_weights[11][40] + inp[41] * layer_1_weights[11][41] + inp[42] * layer_1_weights[11][42] + inp[43] * layer_1_weights[11][43] + inp[44] * layer_1_weights[11][44] + inp[45] * layer_1_weights[11][45] + inp[46] * layer_1_weights[11][46] + inp[47] * layer_1_weights[11][47] + inp[48] * layer_1_weights[11][48] + inp[49] * layer_1_weights[11][49] + inp[50] * layer_1_weights[11][50] + inp[51] * layer_1_weights[11][51] + inp[52] * layer_1_weights[11][52] + inp[53] * layer_1_weights[11][53] + inp[54] * layer_1_weights[11][54] + inp[55] * layer_1_weights[11][55] + inp[56] * layer_1_weights[11][56] + inp[57] * layer_1_weights[11][57] + inp[58] * layer_1_weights[11][58] + inp[59] * layer_1_weights[11][59] + inp[60] * layer_1_weights[11][60] + inp[61] * layer_1_weights[11][61] + inp[62] * layer_1_weights[11][62] + inp[63] * layer_1_weights[11][63] + inp[64] * layer_1_weights[11][64] + inp[65] * layer_1_weights[11][65] + inp[66] * layer_1_weights[11][66] + inp[67] * layer_1_weights[11][67] + inp[68] * layer_1_weights[11][68] + inp[69] * layer_1_weights[11][69] + inp[70] * layer_1_weights[11][70] + inp[71] * layer_1_weights[11][71] + inp[72] * layer_1_weights[11][72] + inp[73] * layer_1_weights[11][73] + inp[74] * layer_1_weights[11][74] + inp[75] * layer_1_weights[11][75] + inp[76] * layer_1_weights[11][76] + inp[77] * layer_1_weights[11][77] + inp[78] * layer_1_weights[11][78] + inp[79] * layer_1_weights[11][79] + inp[80] * layer_1_weights[11][80] + inp[81] * layer_1_weights[11][81] + inp[82] * layer_1_weights[11][82] + inp[83] * layer_1_weights[11][83] + inp[84] * layer_1_weights[11][84] + inp[85] * layer_1_weights[11][85] + inp[86] * layer_1_weights[11][86] + inp[87] * layer_1_weights[11][87] + inp[88] * layer_1_weights[11][88] + inp[89] * layer_1_weights[11][89] + inp[90] * layer_1_weights[11][90] + inp[91] * layer_1_weights[11][91] + inp[92] * layer_1_weights[11][92] + inp[93] * layer_1_weights[11][93] + inp[94] * layer_1_weights[11][94] + inp[95] * layer_1_weights[11][95] + inp[96] * layer_1_weights[11][96] + inp[97] * layer_1_weights[11][97] + inp[98] * layer_1_weights[11][98] + inp[99] * layer_1_weights[11][99] + inp[100] * layer_1_weights[11][100] + inp[101] * layer_1_weights[11][101] + inp[102] * layer_1_weights[11][102] + inp[103] * layer_1_weights[11][103] + inp[104] * layer_1_weights[11][104] + inp[105] * layer_1_weights[11][105] + inp[106] * layer_1_weights[11][106] + inp[107] * layer_1_weights[11][107] + inp[108] * layer_1_weights[11][108] + inp[109] * layer_1_weights[11][109] + inp[110] * layer_1_weights[11][110] + inp[111] * layer_1_weights[11][111] + inp[112] * layer_1_weights[11][112] + inp[113] * layer_1_weights[11][113] + inp[114] * layer_1_weights[11][114] + inp[115] * layer_1_weights[11][115] + inp[116] * layer_1_weights[11][116] + inp[117] * layer_1_weights[11][117] + inp[118] * layer_1_weights[11][118] + inp[119] * layer_1_weights[11][119] + inp[120] * layer_1_weights[11][120] + inp[121] * layer_1_weights[11][121] + inp[122] * layer_1_weights[11][122] + inp[123] * layer_1_weights[11][123] + inp[124] * layer_1_weights[11][124] + inp[125] * layer_1_weights[11][125] + inp[126] * layer_1_weights[11][126] + inp[127] * layer_1_weights[11][127] + inp[128] * layer_1_weights[11][128] + inp[129] * layer_1_weights[11][129] + inp[130] * layer_1_weights[11][130] + inp[131] * layer_1_weights[11][131] + inp[132] * layer_1_weights[11][132] + inp[133] * layer_1_weights[11][133] + inp[134] * layer_1_weights[11][134] + inp[135] * layer_1_weights[11][135] + inp[136] * layer_1_weights[11][136] + inp[137] * layer_1_weights[11][137] + inp[138] * layer_1_weights[11][138] + inp[139] * layer_1_weights[11][139] + inp[140] * layer_1_weights[11][140] + inp[141] * layer_1_weights[11][141] + inp[142] * layer_1_weights[11][142] + inp[143] * layer_1_weights[11][143]);
    assign layer_1_output_12 = relu(layer_1_biases[12] + inp[0] * layer_1_weights[12][0] + inp[1] * layer_1_weights[12][1] + inp[2] * layer_1_weights[12][2] + inp[3] * layer_1_weights[12][3] + inp[4] * layer_1_weights[12][4] + inp[5] * layer_1_weights[12][5] + inp[6] * layer_1_weights[12][6] + inp[7] * layer_1_weights[12][7] + inp[8] * layer_1_weights[12][8] + inp[9] * layer_1_weights[12][9] + inp[10] * layer_1_weights[12][10] + inp[11] * layer_1_weights[12][11] + inp[12] * layer_1_weights[12][12] + inp[13] * layer_1_weights[12][13] + inp[14] * layer_1_weights[12][14] + inp[15] * layer_1_weights[12][15] + inp[16] * layer_1_weights[12][16] + inp[17] * layer_1_weights[12][17] + inp[18] * layer_1_weights[12][18] + inp[19] * layer_1_weights[12][19] + inp[20] * layer_1_weights[12][20] + inp[21] * layer_1_weights[12][21] + inp[22] * layer_1_weights[12][22] + inp[23] * layer_1_weights[12][23] + inp[24] * layer_1_weights[12][24] + inp[25] * layer_1_weights[12][25] + inp[26] * layer_1_weights[12][26] + inp[27] * layer_1_weights[12][27] + inp[28] * layer_1_weights[12][28] + inp[29] * layer_1_weights[12][29] + inp[30] * layer_1_weights[12][30] + inp[31] * layer_1_weights[12][31] + inp[32] * layer_1_weights[12][32] + inp[33] * layer_1_weights[12][33] + inp[34] * layer_1_weights[12][34] + inp[35] * layer_1_weights[12][35] + inp[36] * layer_1_weights[12][36] + inp[37] * layer_1_weights[12][37] + inp[38] * layer_1_weights[12][38] + inp[39] * layer_1_weights[12][39] + inp[40] * layer_1_weights[12][40] + inp[41] * layer_1_weights[12][41] + inp[42] * layer_1_weights[12][42] + inp[43] * layer_1_weights[12][43] + inp[44] * layer_1_weights[12][44] + inp[45] * layer_1_weights[12][45] + inp[46] * layer_1_weights[12][46] + inp[47] * layer_1_weights[12][47] + inp[48] * layer_1_weights[12][48] + inp[49] * layer_1_weights[12][49] + inp[50] * layer_1_weights[12][50] + inp[51] * layer_1_weights[12][51] + inp[52] * layer_1_weights[12][52] + inp[53] * layer_1_weights[12][53] + inp[54] * layer_1_weights[12][54] + inp[55] * layer_1_weights[12][55] + inp[56] * layer_1_weights[12][56] + inp[57] * layer_1_weights[12][57] + inp[58] * layer_1_weights[12][58] + inp[59] * layer_1_weights[12][59] + inp[60] * layer_1_weights[12][60] + inp[61] * layer_1_weights[12][61] + inp[62] * layer_1_weights[12][62] + inp[63] * layer_1_weights[12][63] + inp[64] * layer_1_weights[12][64] + inp[65] * layer_1_weights[12][65] + inp[66] * layer_1_weights[12][66] + inp[67] * layer_1_weights[12][67] + inp[68] * layer_1_weights[12][68] + inp[69] * layer_1_weights[12][69] + inp[70] * layer_1_weights[12][70] + inp[71] * layer_1_weights[12][71] + inp[72] * layer_1_weights[12][72] + inp[73] * layer_1_weights[12][73] + inp[74] * layer_1_weights[12][74] + inp[75] * layer_1_weights[12][75] + inp[76] * layer_1_weights[12][76] + inp[77] * layer_1_weights[12][77] + inp[78] * layer_1_weights[12][78] + inp[79] * layer_1_weights[12][79] + inp[80] * layer_1_weights[12][80] + inp[81] * layer_1_weights[12][81] + inp[82] * layer_1_weights[12][82] + inp[83] * layer_1_weights[12][83] + inp[84] * layer_1_weights[12][84] + inp[85] * layer_1_weights[12][85] + inp[86] * layer_1_weights[12][86] + inp[87] * layer_1_weights[12][87] + inp[88] * layer_1_weights[12][88] + inp[89] * layer_1_weights[12][89] + inp[90] * layer_1_weights[12][90] + inp[91] * layer_1_weights[12][91] + inp[92] * layer_1_weights[12][92] + inp[93] * layer_1_weights[12][93] + inp[94] * layer_1_weights[12][94] + inp[95] * layer_1_weights[12][95] + inp[96] * layer_1_weights[12][96] + inp[97] * layer_1_weights[12][97] + inp[98] * layer_1_weights[12][98] + inp[99] * layer_1_weights[12][99] + inp[100] * layer_1_weights[12][100] + inp[101] * layer_1_weights[12][101] + inp[102] * layer_1_weights[12][102] + inp[103] * layer_1_weights[12][103] + inp[104] * layer_1_weights[12][104] + inp[105] * layer_1_weights[12][105] + inp[106] * layer_1_weights[12][106] + inp[107] * layer_1_weights[12][107] + inp[108] * layer_1_weights[12][108] + inp[109] * layer_1_weights[12][109] + inp[110] * layer_1_weights[12][110] + inp[111] * layer_1_weights[12][111] + inp[112] * layer_1_weights[12][112] + inp[113] * layer_1_weights[12][113] + inp[114] * layer_1_weights[12][114] + inp[115] * layer_1_weights[12][115] + inp[116] * layer_1_weights[12][116] + inp[117] * layer_1_weights[12][117] + inp[118] * layer_1_weights[12][118] + inp[119] * layer_1_weights[12][119] + inp[120] * layer_1_weights[12][120] + inp[121] * layer_1_weights[12][121] + inp[122] * layer_1_weights[12][122] + inp[123] * layer_1_weights[12][123] + inp[124] * layer_1_weights[12][124] + inp[125] * layer_1_weights[12][125] + inp[126] * layer_1_weights[12][126] + inp[127] * layer_1_weights[12][127] + inp[128] * layer_1_weights[12][128] + inp[129] * layer_1_weights[12][129] + inp[130] * layer_1_weights[12][130] + inp[131] * layer_1_weights[12][131] + inp[132] * layer_1_weights[12][132] + inp[133] * layer_1_weights[12][133] + inp[134] * layer_1_weights[12][134] + inp[135] * layer_1_weights[12][135] + inp[136] * layer_1_weights[12][136] + inp[137] * layer_1_weights[12][137] + inp[138] * layer_1_weights[12][138] + inp[139] * layer_1_weights[12][139] + inp[140] * layer_1_weights[12][140] + inp[141] * layer_1_weights[12][141] + inp[142] * layer_1_weights[12][142] + inp[143] * layer_1_weights[12][143]);
    assign layer_1_output_13 = relu(layer_1_biases[13] + inp[0] * layer_1_weights[13][0] + inp[1] * layer_1_weights[13][1] + inp[2] * layer_1_weights[13][2] + inp[3] * layer_1_weights[13][3] + inp[4] * layer_1_weights[13][4] + inp[5] * layer_1_weights[13][5] + inp[6] * layer_1_weights[13][6] + inp[7] * layer_1_weights[13][7] + inp[8] * layer_1_weights[13][8] + inp[9] * layer_1_weights[13][9] + inp[10] * layer_1_weights[13][10] + inp[11] * layer_1_weights[13][11] + inp[12] * layer_1_weights[13][12] + inp[13] * layer_1_weights[13][13] + inp[14] * layer_1_weights[13][14] + inp[15] * layer_1_weights[13][15] + inp[16] * layer_1_weights[13][16] + inp[17] * layer_1_weights[13][17] + inp[18] * layer_1_weights[13][18] + inp[19] * layer_1_weights[13][19] + inp[20] * layer_1_weights[13][20] + inp[21] * layer_1_weights[13][21] + inp[22] * layer_1_weights[13][22] + inp[23] * layer_1_weights[13][23] + inp[24] * layer_1_weights[13][24] + inp[25] * layer_1_weights[13][25] + inp[26] * layer_1_weights[13][26] + inp[27] * layer_1_weights[13][27] + inp[28] * layer_1_weights[13][28] + inp[29] * layer_1_weights[13][29] + inp[30] * layer_1_weights[13][30] + inp[31] * layer_1_weights[13][31] + inp[32] * layer_1_weights[13][32] + inp[33] * layer_1_weights[13][33] + inp[34] * layer_1_weights[13][34] + inp[35] * layer_1_weights[13][35] + inp[36] * layer_1_weights[13][36] + inp[37] * layer_1_weights[13][37] + inp[38] * layer_1_weights[13][38] + inp[39] * layer_1_weights[13][39] + inp[40] * layer_1_weights[13][40] + inp[41] * layer_1_weights[13][41] + inp[42] * layer_1_weights[13][42] + inp[43] * layer_1_weights[13][43] + inp[44] * layer_1_weights[13][44] + inp[45] * layer_1_weights[13][45] + inp[46] * layer_1_weights[13][46] + inp[47] * layer_1_weights[13][47] + inp[48] * layer_1_weights[13][48] + inp[49] * layer_1_weights[13][49] + inp[50] * layer_1_weights[13][50] + inp[51] * layer_1_weights[13][51] + inp[52] * layer_1_weights[13][52] + inp[53] * layer_1_weights[13][53] + inp[54] * layer_1_weights[13][54] + inp[55] * layer_1_weights[13][55] + inp[56] * layer_1_weights[13][56] + inp[57] * layer_1_weights[13][57] + inp[58] * layer_1_weights[13][58] + inp[59] * layer_1_weights[13][59] + inp[60] * layer_1_weights[13][60] + inp[61] * layer_1_weights[13][61] + inp[62] * layer_1_weights[13][62] + inp[63] * layer_1_weights[13][63] + inp[64] * layer_1_weights[13][64] + inp[65] * layer_1_weights[13][65] + inp[66] * layer_1_weights[13][66] + inp[67] * layer_1_weights[13][67] + inp[68] * layer_1_weights[13][68] + inp[69] * layer_1_weights[13][69] + inp[70] * layer_1_weights[13][70] + inp[71] * layer_1_weights[13][71] + inp[72] * layer_1_weights[13][72] + inp[73] * layer_1_weights[13][73] + inp[74] * layer_1_weights[13][74] + inp[75] * layer_1_weights[13][75] + inp[76] * layer_1_weights[13][76] + inp[77] * layer_1_weights[13][77] + inp[78] * layer_1_weights[13][78] + inp[79] * layer_1_weights[13][79] + inp[80] * layer_1_weights[13][80] + inp[81] * layer_1_weights[13][81] + inp[82] * layer_1_weights[13][82] + inp[83] * layer_1_weights[13][83] + inp[84] * layer_1_weights[13][84] + inp[85] * layer_1_weights[13][85] + inp[86] * layer_1_weights[13][86] + inp[87] * layer_1_weights[13][87] + inp[88] * layer_1_weights[13][88] + inp[89] * layer_1_weights[13][89] + inp[90] * layer_1_weights[13][90] + inp[91] * layer_1_weights[13][91] + inp[92] * layer_1_weights[13][92] + inp[93] * layer_1_weights[13][93] + inp[94] * layer_1_weights[13][94] + inp[95] * layer_1_weights[13][95] + inp[96] * layer_1_weights[13][96] + inp[97] * layer_1_weights[13][97] + inp[98] * layer_1_weights[13][98] + inp[99] * layer_1_weights[13][99] + inp[100] * layer_1_weights[13][100] + inp[101] * layer_1_weights[13][101] + inp[102] * layer_1_weights[13][102] + inp[103] * layer_1_weights[13][103] + inp[104] * layer_1_weights[13][104] + inp[105] * layer_1_weights[13][105] + inp[106] * layer_1_weights[13][106] + inp[107] * layer_1_weights[13][107] + inp[108] * layer_1_weights[13][108] + inp[109] * layer_1_weights[13][109] + inp[110] * layer_1_weights[13][110] + inp[111] * layer_1_weights[13][111] + inp[112] * layer_1_weights[13][112] + inp[113] * layer_1_weights[13][113] + inp[114] * layer_1_weights[13][114] + inp[115] * layer_1_weights[13][115] + inp[116] * layer_1_weights[13][116] + inp[117] * layer_1_weights[13][117] + inp[118] * layer_1_weights[13][118] + inp[119] * layer_1_weights[13][119] + inp[120] * layer_1_weights[13][120] + inp[121] * layer_1_weights[13][121] + inp[122] * layer_1_weights[13][122] + inp[123] * layer_1_weights[13][123] + inp[124] * layer_1_weights[13][124] + inp[125] * layer_1_weights[13][125] + inp[126] * layer_1_weights[13][126] + inp[127] * layer_1_weights[13][127] + inp[128] * layer_1_weights[13][128] + inp[129] * layer_1_weights[13][129] + inp[130] * layer_1_weights[13][130] + inp[131] * layer_1_weights[13][131] + inp[132] * layer_1_weights[13][132] + inp[133] * layer_1_weights[13][133] + inp[134] * layer_1_weights[13][134] + inp[135] * layer_1_weights[13][135] + inp[136] * layer_1_weights[13][136] + inp[137] * layer_1_weights[13][137] + inp[138] * layer_1_weights[13][138] + inp[139] * layer_1_weights[13][139] + inp[140] * layer_1_weights[13][140] + inp[141] * layer_1_weights[13][141] + inp[142] * layer_1_weights[13][142] + inp[143] * layer_1_weights[13][143]);
    assign layer_1_output_14 = relu(layer_1_biases[14] + inp[0] * layer_1_weights[14][0] + inp[1] * layer_1_weights[14][1] + inp[2] * layer_1_weights[14][2] + inp[3] * layer_1_weights[14][3] + inp[4] * layer_1_weights[14][4] + inp[5] * layer_1_weights[14][5] + inp[6] * layer_1_weights[14][6] + inp[7] * layer_1_weights[14][7] + inp[8] * layer_1_weights[14][8] + inp[9] * layer_1_weights[14][9] + inp[10] * layer_1_weights[14][10] + inp[11] * layer_1_weights[14][11] + inp[12] * layer_1_weights[14][12] + inp[13] * layer_1_weights[14][13] + inp[14] * layer_1_weights[14][14] + inp[15] * layer_1_weights[14][15] + inp[16] * layer_1_weights[14][16] + inp[17] * layer_1_weights[14][17] + inp[18] * layer_1_weights[14][18] + inp[19] * layer_1_weights[14][19] + inp[20] * layer_1_weights[14][20] + inp[21] * layer_1_weights[14][21] + inp[22] * layer_1_weights[14][22] + inp[23] * layer_1_weights[14][23] + inp[24] * layer_1_weights[14][24] + inp[25] * layer_1_weights[14][25] + inp[26] * layer_1_weights[14][26] + inp[27] * layer_1_weights[14][27] + inp[28] * layer_1_weights[14][28] + inp[29] * layer_1_weights[14][29] + inp[30] * layer_1_weights[14][30] + inp[31] * layer_1_weights[14][31] + inp[32] * layer_1_weights[14][32] + inp[33] * layer_1_weights[14][33] + inp[34] * layer_1_weights[14][34] + inp[35] * layer_1_weights[14][35] + inp[36] * layer_1_weights[14][36] + inp[37] * layer_1_weights[14][37] + inp[38] * layer_1_weights[14][38] + inp[39] * layer_1_weights[14][39] + inp[40] * layer_1_weights[14][40] + inp[41] * layer_1_weights[14][41] + inp[42] * layer_1_weights[14][42] + inp[43] * layer_1_weights[14][43] + inp[44] * layer_1_weights[14][44] + inp[45] * layer_1_weights[14][45] + inp[46] * layer_1_weights[14][46] + inp[47] * layer_1_weights[14][47] + inp[48] * layer_1_weights[14][48] + inp[49] * layer_1_weights[14][49] + inp[50] * layer_1_weights[14][50] + inp[51] * layer_1_weights[14][51] + inp[52] * layer_1_weights[14][52] + inp[53] * layer_1_weights[14][53] + inp[54] * layer_1_weights[14][54] + inp[55] * layer_1_weights[14][55] + inp[56] * layer_1_weights[14][56] + inp[57] * layer_1_weights[14][57] + inp[58] * layer_1_weights[14][58] + inp[59] * layer_1_weights[14][59] + inp[60] * layer_1_weights[14][60] + inp[61] * layer_1_weights[14][61] + inp[62] * layer_1_weights[14][62] + inp[63] * layer_1_weights[14][63] + inp[64] * layer_1_weights[14][64] + inp[65] * layer_1_weights[14][65] + inp[66] * layer_1_weights[14][66] + inp[67] * layer_1_weights[14][67] + inp[68] * layer_1_weights[14][68] + inp[69] * layer_1_weights[14][69] + inp[70] * layer_1_weights[14][70] + inp[71] * layer_1_weights[14][71] + inp[72] * layer_1_weights[14][72] + inp[73] * layer_1_weights[14][73] + inp[74] * layer_1_weights[14][74] + inp[75] * layer_1_weights[14][75] + inp[76] * layer_1_weights[14][76] + inp[77] * layer_1_weights[14][77] + inp[78] * layer_1_weights[14][78] + inp[79] * layer_1_weights[14][79] + inp[80] * layer_1_weights[14][80] + inp[81] * layer_1_weights[14][81] + inp[82] * layer_1_weights[14][82] + inp[83] * layer_1_weights[14][83] + inp[84] * layer_1_weights[14][84] + inp[85] * layer_1_weights[14][85] + inp[86] * layer_1_weights[14][86] + inp[87] * layer_1_weights[14][87] + inp[88] * layer_1_weights[14][88] + inp[89] * layer_1_weights[14][89] + inp[90] * layer_1_weights[14][90] + inp[91] * layer_1_weights[14][91] + inp[92] * layer_1_weights[14][92] + inp[93] * layer_1_weights[14][93] + inp[94] * layer_1_weights[14][94] + inp[95] * layer_1_weights[14][95] + inp[96] * layer_1_weights[14][96] + inp[97] * layer_1_weights[14][97] + inp[98] * layer_1_weights[14][98] + inp[99] * layer_1_weights[14][99] + inp[100] * layer_1_weights[14][100] + inp[101] * layer_1_weights[14][101] + inp[102] * layer_1_weights[14][102] + inp[103] * layer_1_weights[14][103] + inp[104] * layer_1_weights[14][104] + inp[105] * layer_1_weights[14][105] + inp[106] * layer_1_weights[14][106] + inp[107] * layer_1_weights[14][107] + inp[108] * layer_1_weights[14][108] + inp[109] * layer_1_weights[14][109] + inp[110] * layer_1_weights[14][110] + inp[111] * layer_1_weights[14][111] + inp[112] * layer_1_weights[14][112] + inp[113] * layer_1_weights[14][113] + inp[114] * layer_1_weights[14][114] + inp[115] * layer_1_weights[14][115] + inp[116] * layer_1_weights[14][116] + inp[117] * layer_1_weights[14][117] + inp[118] * layer_1_weights[14][118] + inp[119] * layer_1_weights[14][119] + inp[120] * layer_1_weights[14][120] + inp[121] * layer_1_weights[14][121] + inp[122] * layer_1_weights[14][122] + inp[123] * layer_1_weights[14][123] + inp[124] * layer_1_weights[14][124] + inp[125] * layer_1_weights[14][125] + inp[126] * layer_1_weights[14][126] + inp[127] * layer_1_weights[14][127] + inp[128] * layer_1_weights[14][128] + inp[129] * layer_1_weights[14][129] + inp[130] * layer_1_weights[14][130] + inp[131] * layer_1_weights[14][131] + inp[132] * layer_1_weights[14][132] + inp[133] * layer_1_weights[14][133] + inp[134] * layer_1_weights[14][134] + inp[135] * layer_1_weights[14][135] + inp[136] * layer_1_weights[14][136] + inp[137] * layer_1_weights[14][137] + inp[138] * layer_1_weights[14][138] + inp[139] * layer_1_weights[14][139] + inp[140] * layer_1_weights[14][140] + inp[141] * layer_1_weights[14][141] + inp[142] * layer_1_weights[14][142] + inp[143] * layer_1_weights[14][143]);
    assign layer_1_output_15 = relu(layer_1_biases[15] + inp[0] * layer_1_weights[15][0] + inp[1] * layer_1_weights[15][1] + inp[2] * layer_1_weights[15][2] + inp[3] * layer_1_weights[15][3] + inp[4] * layer_1_weights[15][4] + inp[5] * layer_1_weights[15][5] + inp[6] * layer_1_weights[15][6] + inp[7] * layer_1_weights[15][7] + inp[8] * layer_1_weights[15][8] + inp[9] * layer_1_weights[15][9] + inp[10] * layer_1_weights[15][10] + inp[11] * layer_1_weights[15][11] + inp[12] * layer_1_weights[15][12] + inp[13] * layer_1_weights[15][13] + inp[14] * layer_1_weights[15][14] + inp[15] * layer_1_weights[15][15] + inp[16] * layer_1_weights[15][16] + inp[17] * layer_1_weights[15][17] + inp[18] * layer_1_weights[15][18] + inp[19] * layer_1_weights[15][19] + inp[20] * layer_1_weights[15][20] + inp[21] * layer_1_weights[15][21] + inp[22] * layer_1_weights[15][22] + inp[23] * layer_1_weights[15][23] + inp[24] * layer_1_weights[15][24] + inp[25] * layer_1_weights[15][25] + inp[26] * layer_1_weights[15][26] + inp[27] * layer_1_weights[15][27] + inp[28] * layer_1_weights[15][28] + inp[29] * layer_1_weights[15][29] + inp[30] * layer_1_weights[15][30] + inp[31] * layer_1_weights[15][31] + inp[32] * layer_1_weights[15][32] + inp[33] * layer_1_weights[15][33] + inp[34] * layer_1_weights[15][34] + inp[35] * layer_1_weights[15][35] + inp[36] * layer_1_weights[15][36] + inp[37] * layer_1_weights[15][37] + inp[38] * layer_1_weights[15][38] + inp[39] * layer_1_weights[15][39] + inp[40] * layer_1_weights[15][40] + inp[41] * layer_1_weights[15][41] + inp[42] * layer_1_weights[15][42] + inp[43] * layer_1_weights[15][43] + inp[44] * layer_1_weights[15][44] + inp[45] * layer_1_weights[15][45] + inp[46] * layer_1_weights[15][46] + inp[47] * layer_1_weights[15][47] + inp[48] * layer_1_weights[15][48] + inp[49] * layer_1_weights[15][49] + inp[50] * layer_1_weights[15][50] + inp[51] * layer_1_weights[15][51] + inp[52] * layer_1_weights[15][52] + inp[53] * layer_1_weights[15][53] + inp[54] * layer_1_weights[15][54] + inp[55] * layer_1_weights[15][55] + inp[56] * layer_1_weights[15][56] + inp[57] * layer_1_weights[15][57] + inp[58] * layer_1_weights[15][58] + inp[59] * layer_1_weights[15][59] + inp[60] * layer_1_weights[15][60] + inp[61] * layer_1_weights[15][61] + inp[62] * layer_1_weights[15][62] + inp[63] * layer_1_weights[15][63] + inp[64] * layer_1_weights[15][64] + inp[65] * layer_1_weights[15][65] + inp[66] * layer_1_weights[15][66] + inp[67] * layer_1_weights[15][67] + inp[68] * layer_1_weights[15][68] + inp[69] * layer_1_weights[15][69] + inp[70] * layer_1_weights[15][70] + inp[71] * layer_1_weights[15][71] + inp[72] * layer_1_weights[15][72] + inp[73] * layer_1_weights[15][73] + inp[74] * layer_1_weights[15][74] + inp[75] * layer_1_weights[15][75] + inp[76] * layer_1_weights[15][76] + inp[77] * layer_1_weights[15][77] + inp[78] * layer_1_weights[15][78] + inp[79] * layer_1_weights[15][79] + inp[80] * layer_1_weights[15][80] + inp[81] * layer_1_weights[15][81] + inp[82] * layer_1_weights[15][82] + inp[83] * layer_1_weights[15][83] + inp[84] * layer_1_weights[15][84] + inp[85] * layer_1_weights[15][85] + inp[86] * layer_1_weights[15][86] + inp[87] * layer_1_weights[15][87] + inp[88] * layer_1_weights[15][88] + inp[89] * layer_1_weights[15][89] + inp[90] * layer_1_weights[15][90] + inp[91] * layer_1_weights[15][91] + inp[92] * layer_1_weights[15][92] + inp[93] * layer_1_weights[15][93] + inp[94] * layer_1_weights[15][94] + inp[95] * layer_1_weights[15][95] + inp[96] * layer_1_weights[15][96] + inp[97] * layer_1_weights[15][97] + inp[98] * layer_1_weights[15][98] + inp[99] * layer_1_weights[15][99] + inp[100] * layer_1_weights[15][100] + inp[101] * layer_1_weights[15][101] + inp[102] * layer_1_weights[15][102] + inp[103] * layer_1_weights[15][103] + inp[104] * layer_1_weights[15][104] + inp[105] * layer_1_weights[15][105] + inp[106] * layer_1_weights[15][106] + inp[107] * layer_1_weights[15][107] + inp[108] * layer_1_weights[15][108] + inp[109] * layer_1_weights[15][109] + inp[110] * layer_1_weights[15][110] + inp[111] * layer_1_weights[15][111] + inp[112] * layer_1_weights[15][112] + inp[113] * layer_1_weights[15][113] + inp[114] * layer_1_weights[15][114] + inp[115] * layer_1_weights[15][115] + inp[116] * layer_1_weights[15][116] + inp[117] * layer_1_weights[15][117] + inp[118] * layer_1_weights[15][118] + inp[119] * layer_1_weights[15][119] + inp[120] * layer_1_weights[15][120] + inp[121] * layer_1_weights[15][121] + inp[122] * layer_1_weights[15][122] + inp[123] * layer_1_weights[15][123] + inp[124] * layer_1_weights[15][124] + inp[125] * layer_1_weights[15][125] + inp[126] * layer_1_weights[15][126] + inp[127] * layer_1_weights[15][127] + inp[128] * layer_1_weights[15][128] + inp[129] * layer_1_weights[15][129] + inp[130] * layer_1_weights[15][130] + inp[131] * layer_1_weights[15][131] + inp[132] * layer_1_weights[15][132] + inp[133] * layer_1_weights[15][133] + inp[134] * layer_1_weights[15][134] + inp[135] * layer_1_weights[15][135] + inp[136] * layer_1_weights[15][136] + inp[137] * layer_1_weights[15][137] + inp[138] * layer_1_weights[15][138] + inp[139] * layer_1_weights[15][139] + inp[140] * layer_1_weights[15][140] + inp[141] * layer_1_weights[15][141] + inp[142] * layer_1_weights[15][142] + inp[143] * layer_1_weights[15][143]);
    assign layer_1_output_16 = relu(layer_1_biases[16] + inp[0] * layer_1_weights[16][0] + inp[1] * layer_1_weights[16][1] + inp[2] * layer_1_weights[16][2] + inp[3] * layer_1_weights[16][3] + inp[4] * layer_1_weights[16][4] + inp[5] * layer_1_weights[16][5] + inp[6] * layer_1_weights[16][6] + inp[7] * layer_1_weights[16][7] + inp[8] * layer_1_weights[16][8] + inp[9] * layer_1_weights[16][9] + inp[10] * layer_1_weights[16][10] + inp[11] * layer_1_weights[16][11] + inp[12] * layer_1_weights[16][12] + inp[13] * layer_1_weights[16][13] + inp[14] * layer_1_weights[16][14] + inp[15] * layer_1_weights[16][15] + inp[16] * layer_1_weights[16][16] + inp[17] * layer_1_weights[16][17] + inp[18] * layer_1_weights[16][18] + inp[19] * layer_1_weights[16][19] + inp[20] * layer_1_weights[16][20] + inp[21] * layer_1_weights[16][21] + inp[22] * layer_1_weights[16][22] + inp[23] * layer_1_weights[16][23] + inp[24] * layer_1_weights[16][24] + inp[25] * layer_1_weights[16][25] + inp[26] * layer_1_weights[16][26] + inp[27] * layer_1_weights[16][27] + inp[28] * layer_1_weights[16][28] + inp[29] * layer_1_weights[16][29] + inp[30] * layer_1_weights[16][30] + inp[31] * layer_1_weights[16][31] + inp[32] * layer_1_weights[16][32] + inp[33] * layer_1_weights[16][33] + inp[34] * layer_1_weights[16][34] + inp[35] * layer_1_weights[16][35] + inp[36] * layer_1_weights[16][36] + inp[37] * layer_1_weights[16][37] + inp[38] * layer_1_weights[16][38] + inp[39] * layer_1_weights[16][39] + inp[40] * layer_1_weights[16][40] + inp[41] * layer_1_weights[16][41] + inp[42] * layer_1_weights[16][42] + inp[43] * layer_1_weights[16][43] + inp[44] * layer_1_weights[16][44] + inp[45] * layer_1_weights[16][45] + inp[46] * layer_1_weights[16][46] + inp[47] * layer_1_weights[16][47] + inp[48] * layer_1_weights[16][48] + inp[49] * layer_1_weights[16][49] + inp[50] * layer_1_weights[16][50] + inp[51] * layer_1_weights[16][51] + inp[52] * layer_1_weights[16][52] + inp[53] * layer_1_weights[16][53] + inp[54] * layer_1_weights[16][54] + inp[55] * layer_1_weights[16][55] + inp[56] * layer_1_weights[16][56] + inp[57] * layer_1_weights[16][57] + inp[58] * layer_1_weights[16][58] + inp[59] * layer_1_weights[16][59] + inp[60] * layer_1_weights[16][60] + inp[61] * layer_1_weights[16][61] + inp[62] * layer_1_weights[16][62] + inp[63] * layer_1_weights[16][63] + inp[64] * layer_1_weights[16][64] + inp[65] * layer_1_weights[16][65] + inp[66] * layer_1_weights[16][66] + inp[67] * layer_1_weights[16][67] + inp[68] * layer_1_weights[16][68] + inp[69] * layer_1_weights[16][69] + inp[70] * layer_1_weights[16][70] + inp[71] * layer_1_weights[16][71] + inp[72] * layer_1_weights[16][72] + inp[73] * layer_1_weights[16][73] + inp[74] * layer_1_weights[16][74] + inp[75] * layer_1_weights[16][75] + inp[76] * layer_1_weights[16][76] + inp[77] * layer_1_weights[16][77] + inp[78] * layer_1_weights[16][78] + inp[79] * layer_1_weights[16][79] + inp[80] * layer_1_weights[16][80] + inp[81] * layer_1_weights[16][81] + inp[82] * layer_1_weights[16][82] + inp[83] * layer_1_weights[16][83] + inp[84] * layer_1_weights[16][84] + inp[85] * layer_1_weights[16][85] + inp[86] * layer_1_weights[16][86] + inp[87] * layer_1_weights[16][87] + inp[88] * layer_1_weights[16][88] + inp[89] * layer_1_weights[16][89] + inp[90] * layer_1_weights[16][90] + inp[91] * layer_1_weights[16][91] + inp[92] * layer_1_weights[16][92] + inp[93] * layer_1_weights[16][93] + inp[94] * layer_1_weights[16][94] + inp[95] * layer_1_weights[16][95] + inp[96] * layer_1_weights[16][96] + inp[97] * layer_1_weights[16][97] + inp[98] * layer_1_weights[16][98] + inp[99] * layer_1_weights[16][99] + inp[100] * layer_1_weights[16][100] + inp[101] * layer_1_weights[16][101] + inp[102] * layer_1_weights[16][102] + inp[103] * layer_1_weights[16][103] + inp[104] * layer_1_weights[16][104] + inp[105] * layer_1_weights[16][105] + inp[106] * layer_1_weights[16][106] + inp[107] * layer_1_weights[16][107] + inp[108] * layer_1_weights[16][108] + inp[109] * layer_1_weights[16][109] + inp[110] * layer_1_weights[16][110] + inp[111] * layer_1_weights[16][111] + inp[112] * layer_1_weights[16][112] + inp[113] * layer_1_weights[16][113] + inp[114] * layer_1_weights[16][114] + inp[115] * layer_1_weights[16][115] + inp[116] * layer_1_weights[16][116] + inp[117] * layer_1_weights[16][117] + inp[118] * layer_1_weights[16][118] + inp[119] * layer_1_weights[16][119] + inp[120] * layer_1_weights[16][120] + inp[121] * layer_1_weights[16][121] + inp[122] * layer_1_weights[16][122] + inp[123] * layer_1_weights[16][123] + inp[124] * layer_1_weights[16][124] + inp[125] * layer_1_weights[16][125] + inp[126] * layer_1_weights[16][126] + inp[127] * layer_1_weights[16][127] + inp[128] * layer_1_weights[16][128] + inp[129] * layer_1_weights[16][129] + inp[130] * layer_1_weights[16][130] + inp[131] * layer_1_weights[16][131] + inp[132] * layer_1_weights[16][132] + inp[133] * layer_1_weights[16][133] + inp[134] * layer_1_weights[16][134] + inp[135] * layer_1_weights[16][135] + inp[136] * layer_1_weights[16][136] + inp[137] * layer_1_weights[16][137] + inp[138] * layer_1_weights[16][138] + inp[139] * layer_1_weights[16][139] + inp[140] * layer_1_weights[16][140] + inp[141] * layer_1_weights[16][141] + inp[142] * layer_1_weights[16][142] + inp[143] * layer_1_weights[16][143]);
    assign layer_1_output_17 = relu(layer_1_biases[17] + inp[0] * layer_1_weights[17][0] + inp[1] * layer_1_weights[17][1] + inp[2] * layer_1_weights[17][2] + inp[3] * layer_1_weights[17][3] + inp[4] * layer_1_weights[17][4] + inp[5] * layer_1_weights[17][5] + inp[6] * layer_1_weights[17][6] + inp[7] * layer_1_weights[17][7] + inp[8] * layer_1_weights[17][8] + inp[9] * layer_1_weights[17][9] + inp[10] * layer_1_weights[17][10] + inp[11] * layer_1_weights[17][11] + inp[12] * layer_1_weights[17][12] + inp[13] * layer_1_weights[17][13] + inp[14] * layer_1_weights[17][14] + inp[15] * layer_1_weights[17][15] + inp[16] * layer_1_weights[17][16] + inp[17] * layer_1_weights[17][17] + inp[18] * layer_1_weights[17][18] + inp[19] * layer_1_weights[17][19] + inp[20] * layer_1_weights[17][20] + inp[21] * layer_1_weights[17][21] + inp[22] * layer_1_weights[17][22] + inp[23] * layer_1_weights[17][23] + inp[24] * layer_1_weights[17][24] + inp[25] * layer_1_weights[17][25] + inp[26] * layer_1_weights[17][26] + inp[27] * layer_1_weights[17][27] + inp[28] * layer_1_weights[17][28] + inp[29] * layer_1_weights[17][29] + inp[30] * layer_1_weights[17][30] + inp[31] * layer_1_weights[17][31] + inp[32] * layer_1_weights[17][32] + inp[33] * layer_1_weights[17][33] + inp[34] * layer_1_weights[17][34] + inp[35] * layer_1_weights[17][35] + inp[36] * layer_1_weights[17][36] + inp[37] * layer_1_weights[17][37] + inp[38] * layer_1_weights[17][38] + inp[39] * layer_1_weights[17][39] + inp[40] * layer_1_weights[17][40] + inp[41] * layer_1_weights[17][41] + inp[42] * layer_1_weights[17][42] + inp[43] * layer_1_weights[17][43] + inp[44] * layer_1_weights[17][44] + inp[45] * layer_1_weights[17][45] + inp[46] * layer_1_weights[17][46] + inp[47] * layer_1_weights[17][47] + inp[48] * layer_1_weights[17][48] + inp[49] * layer_1_weights[17][49] + inp[50] * layer_1_weights[17][50] + inp[51] * layer_1_weights[17][51] + inp[52] * layer_1_weights[17][52] + inp[53] * layer_1_weights[17][53] + inp[54] * layer_1_weights[17][54] + inp[55] * layer_1_weights[17][55] + inp[56] * layer_1_weights[17][56] + inp[57] * layer_1_weights[17][57] + inp[58] * layer_1_weights[17][58] + inp[59] * layer_1_weights[17][59] + inp[60] * layer_1_weights[17][60] + inp[61] * layer_1_weights[17][61] + inp[62] * layer_1_weights[17][62] + inp[63] * layer_1_weights[17][63] + inp[64] * layer_1_weights[17][64] + inp[65] * layer_1_weights[17][65] + inp[66] * layer_1_weights[17][66] + inp[67] * layer_1_weights[17][67] + inp[68] * layer_1_weights[17][68] + inp[69] * layer_1_weights[17][69] + inp[70] * layer_1_weights[17][70] + inp[71] * layer_1_weights[17][71] + inp[72] * layer_1_weights[17][72] + inp[73] * layer_1_weights[17][73] + inp[74] * layer_1_weights[17][74] + inp[75] * layer_1_weights[17][75] + inp[76] * layer_1_weights[17][76] + inp[77] * layer_1_weights[17][77] + inp[78] * layer_1_weights[17][78] + inp[79] * layer_1_weights[17][79] + inp[80] * layer_1_weights[17][80] + inp[81] * layer_1_weights[17][81] + inp[82] * layer_1_weights[17][82] + inp[83] * layer_1_weights[17][83] + inp[84] * layer_1_weights[17][84] + inp[85] * layer_1_weights[17][85] + inp[86] * layer_1_weights[17][86] + inp[87] * layer_1_weights[17][87] + inp[88] * layer_1_weights[17][88] + inp[89] * layer_1_weights[17][89] + inp[90] * layer_1_weights[17][90] + inp[91] * layer_1_weights[17][91] + inp[92] * layer_1_weights[17][92] + inp[93] * layer_1_weights[17][93] + inp[94] * layer_1_weights[17][94] + inp[95] * layer_1_weights[17][95] + inp[96] * layer_1_weights[17][96] + inp[97] * layer_1_weights[17][97] + inp[98] * layer_1_weights[17][98] + inp[99] * layer_1_weights[17][99] + inp[100] * layer_1_weights[17][100] + inp[101] * layer_1_weights[17][101] + inp[102] * layer_1_weights[17][102] + inp[103] * layer_1_weights[17][103] + inp[104] * layer_1_weights[17][104] + inp[105] * layer_1_weights[17][105] + inp[106] * layer_1_weights[17][106] + inp[107] * layer_1_weights[17][107] + inp[108] * layer_1_weights[17][108] + inp[109] * layer_1_weights[17][109] + inp[110] * layer_1_weights[17][110] + inp[111] * layer_1_weights[17][111] + inp[112] * layer_1_weights[17][112] + inp[113] * layer_1_weights[17][113] + inp[114] * layer_1_weights[17][114] + inp[115] * layer_1_weights[17][115] + inp[116] * layer_1_weights[17][116] + inp[117] * layer_1_weights[17][117] + inp[118] * layer_1_weights[17][118] + inp[119] * layer_1_weights[17][119] + inp[120] * layer_1_weights[17][120] + inp[121] * layer_1_weights[17][121] + inp[122] * layer_1_weights[17][122] + inp[123] * layer_1_weights[17][123] + inp[124] * layer_1_weights[17][124] + inp[125] * layer_1_weights[17][125] + inp[126] * layer_1_weights[17][126] + inp[127] * layer_1_weights[17][127] + inp[128] * layer_1_weights[17][128] + inp[129] * layer_1_weights[17][129] + inp[130] * layer_1_weights[17][130] + inp[131] * layer_1_weights[17][131] + inp[132] * layer_1_weights[17][132] + inp[133] * layer_1_weights[17][133] + inp[134] * layer_1_weights[17][134] + inp[135] * layer_1_weights[17][135] + inp[136] * layer_1_weights[17][136] + inp[137] * layer_1_weights[17][137] + inp[138] * layer_1_weights[17][138] + inp[139] * layer_1_weights[17][139] + inp[140] * layer_1_weights[17][140] + inp[141] * layer_1_weights[17][141] + inp[142] * layer_1_weights[17][142] + inp[143] * layer_1_weights[17][143]);
    assign layer_1_output_18 = relu(layer_1_biases[18] + inp[0] * layer_1_weights[18][0] + inp[1] * layer_1_weights[18][1] + inp[2] * layer_1_weights[18][2] + inp[3] * layer_1_weights[18][3] + inp[4] * layer_1_weights[18][4] + inp[5] * layer_1_weights[18][5] + inp[6] * layer_1_weights[18][6] + inp[7] * layer_1_weights[18][7] + inp[8] * layer_1_weights[18][8] + inp[9] * layer_1_weights[18][9] + inp[10] * layer_1_weights[18][10] + inp[11] * layer_1_weights[18][11] + inp[12] * layer_1_weights[18][12] + inp[13] * layer_1_weights[18][13] + inp[14] * layer_1_weights[18][14] + inp[15] * layer_1_weights[18][15] + inp[16] * layer_1_weights[18][16] + inp[17] * layer_1_weights[18][17] + inp[18] * layer_1_weights[18][18] + inp[19] * layer_1_weights[18][19] + inp[20] * layer_1_weights[18][20] + inp[21] * layer_1_weights[18][21] + inp[22] * layer_1_weights[18][22] + inp[23] * layer_1_weights[18][23] + inp[24] * layer_1_weights[18][24] + inp[25] * layer_1_weights[18][25] + inp[26] * layer_1_weights[18][26] + inp[27] * layer_1_weights[18][27] + inp[28] * layer_1_weights[18][28] + inp[29] * layer_1_weights[18][29] + inp[30] * layer_1_weights[18][30] + inp[31] * layer_1_weights[18][31] + inp[32] * layer_1_weights[18][32] + inp[33] * layer_1_weights[18][33] + inp[34] * layer_1_weights[18][34] + inp[35] * layer_1_weights[18][35] + inp[36] * layer_1_weights[18][36] + inp[37] * layer_1_weights[18][37] + inp[38] * layer_1_weights[18][38] + inp[39] * layer_1_weights[18][39] + inp[40] * layer_1_weights[18][40] + inp[41] * layer_1_weights[18][41] + inp[42] * layer_1_weights[18][42] + inp[43] * layer_1_weights[18][43] + inp[44] * layer_1_weights[18][44] + inp[45] * layer_1_weights[18][45] + inp[46] * layer_1_weights[18][46] + inp[47] * layer_1_weights[18][47] + inp[48] * layer_1_weights[18][48] + inp[49] * layer_1_weights[18][49] + inp[50] * layer_1_weights[18][50] + inp[51] * layer_1_weights[18][51] + inp[52] * layer_1_weights[18][52] + inp[53] * layer_1_weights[18][53] + inp[54] * layer_1_weights[18][54] + inp[55] * layer_1_weights[18][55] + inp[56] * layer_1_weights[18][56] + inp[57] * layer_1_weights[18][57] + inp[58] * layer_1_weights[18][58] + inp[59] * layer_1_weights[18][59] + inp[60] * layer_1_weights[18][60] + inp[61] * layer_1_weights[18][61] + inp[62] * layer_1_weights[18][62] + inp[63] * layer_1_weights[18][63] + inp[64] * layer_1_weights[18][64] + inp[65] * layer_1_weights[18][65] + inp[66] * layer_1_weights[18][66] + inp[67] * layer_1_weights[18][67] + inp[68] * layer_1_weights[18][68] + inp[69] * layer_1_weights[18][69] + inp[70] * layer_1_weights[18][70] + inp[71] * layer_1_weights[18][71] + inp[72] * layer_1_weights[18][72] + inp[73] * layer_1_weights[18][73] + inp[74] * layer_1_weights[18][74] + inp[75] * layer_1_weights[18][75] + inp[76] * layer_1_weights[18][76] + inp[77] * layer_1_weights[18][77] + inp[78] * layer_1_weights[18][78] + inp[79] * layer_1_weights[18][79] + inp[80] * layer_1_weights[18][80] + inp[81] * layer_1_weights[18][81] + inp[82] * layer_1_weights[18][82] + inp[83] * layer_1_weights[18][83] + inp[84] * layer_1_weights[18][84] + inp[85] * layer_1_weights[18][85] + inp[86] * layer_1_weights[18][86] + inp[87] * layer_1_weights[18][87] + inp[88] * layer_1_weights[18][88] + inp[89] * layer_1_weights[18][89] + inp[90] * layer_1_weights[18][90] + inp[91] * layer_1_weights[18][91] + inp[92] * layer_1_weights[18][92] + inp[93] * layer_1_weights[18][93] + inp[94] * layer_1_weights[18][94] + inp[95] * layer_1_weights[18][95] + inp[96] * layer_1_weights[18][96] + inp[97] * layer_1_weights[18][97] + inp[98] * layer_1_weights[18][98] + inp[99] * layer_1_weights[18][99] + inp[100] * layer_1_weights[18][100] + inp[101] * layer_1_weights[18][101] + inp[102] * layer_1_weights[18][102] + inp[103] * layer_1_weights[18][103] + inp[104] * layer_1_weights[18][104] + inp[105] * layer_1_weights[18][105] + inp[106] * layer_1_weights[18][106] + inp[107] * layer_1_weights[18][107] + inp[108] * layer_1_weights[18][108] + inp[109] * layer_1_weights[18][109] + inp[110] * layer_1_weights[18][110] + inp[111] * layer_1_weights[18][111] + inp[112] * layer_1_weights[18][112] + inp[113] * layer_1_weights[18][113] + inp[114] * layer_1_weights[18][114] + inp[115] * layer_1_weights[18][115] + inp[116] * layer_1_weights[18][116] + inp[117] * layer_1_weights[18][117] + inp[118] * layer_1_weights[18][118] + inp[119] * layer_1_weights[18][119] + inp[120] * layer_1_weights[18][120] + inp[121] * layer_1_weights[18][121] + inp[122] * layer_1_weights[18][122] + inp[123] * layer_1_weights[18][123] + inp[124] * layer_1_weights[18][124] + inp[125] * layer_1_weights[18][125] + inp[126] * layer_1_weights[18][126] + inp[127] * layer_1_weights[18][127] + inp[128] * layer_1_weights[18][128] + inp[129] * layer_1_weights[18][129] + inp[130] * layer_1_weights[18][130] + inp[131] * layer_1_weights[18][131] + inp[132] * layer_1_weights[18][132] + inp[133] * layer_1_weights[18][133] + inp[134] * layer_1_weights[18][134] + inp[135] * layer_1_weights[18][135] + inp[136] * layer_1_weights[18][136] + inp[137] * layer_1_weights[18][137] + inp[138] * layer_1_weights[18][138] + inp[139] * layer_1_weights[18][139] + inp[140] * layer_1_weights[18][140] + inp[141] * layer_1_weights[18][141] + inp[142] * layer_1_weights[18][142] + inp[143] * layer_1_weights[18][143]);
    assign layer_1_output_19 = relu(layer_1_biases[19] + inp[0] * layer_1_weights[19][0] + inp[1] * layer_1_weights[19][1] + inp[2] * layer_1_weights[19][2] + inp[3] * layer_1_weights[19][3] + inp[4] * layer_1_weights[19][4] + inp[5] * layer_1_weights[19][5] + inp[6] * layer_1_weights[19][6] + inp[7] * layer_1_weights[19][7] + inp[8] * layer_1_weights[19][8] + inp[9] * layer_1_weights[19][9] + inp[10] * layer_1_weights[19][10] + inp[11] * layer_1_weights[19][11] + inp[12] * layer_1_weights[19][12] + inp[13] * layer_1_weights[19][13] + inp[14] * layer_1_weights[19][14] + inp[15] * layer_1_weights[19][15] + inp[16] * layer_1_weights[19][16] + inp[17] * layer_1_weights[19][17] + inp[18] * layer_1_weights[19][18] + inp[19] * layer_1_weights[19][19] + inp[20] * layer_1_weights[19][20] + inp[21] * layer_1_weights[19][21] + inp[22] * layer_1_weights[19][22] + inp[23] * layer_1_weights[19][23] + inp[24] * layer_1_weights[19][24] + inp[25] * layer_1_weights[19][25] + inp[26] * layer_1_weights[19][26] + inp[27] * layer_1_weights[19][27] + inp[28] * layer_1_weights[19][28] + inp[29] * layer_1_weights[19][29] + inp[30] * layer_1_weights[19][30] + inp[31] * layer_1_weights[19][31] + inp[32] * layer_1_weights[19][32] + inp[33] * layer_1_weights[19][33] + inp[34] * layer_1_weights[19][34] + inp[35] * layer_1_weights[19][35] + inp[36] * layer_1_weights[19][36] + inp[37] * layer_1_weights[19][37] + inp[38] * layer_1_weights[19][38] + inp[39] * layer_1_weights[19][39] + inp[40] * layer_1_weights[19][40] + inp[41] * layer_1_weights[19][41] + inp[42] * layer_1_weights[19][42] + inp[43] * layer_1_weights[19][43] + inp[44] * layer_1_weights[19][44] + inp[45] * layer_1_weights[19][45] + inp[46] * layer_1_weights[19][46] + inp[47] * layer_1_weights[19][47] + inp[48] * layer_1_weights[19][48] + inp[49] * layer_1_weights[19][49] + inp[50] * layer_1_weights[19][50] + inp[51] * layer_1_weights[19][51] + inp[52] * layer_1_weights[19][52] + inp[53] * layer_1_weights[19][53] + inp[54] * layer_1_weights[19][54] + inp[55] * layer_1_weights[19][55] + inp[56] * layer_1_weights[19][56] + inp[57] * layer_1_weights[19][57] + inp[58] * layer_1_weights[19][58] + inp[59] * layer_1_weights[19][59] + inp[60] * layer_1_weights[19][60] + inp[61] * layer_1_weights[19][61] + inp[62] * layer_1_weights[19][62] + inp[63] * layer_1_weights[19][63] + inp[64] * layer_1_weights[19][64] + inp[65] * layer_1_weights[19][65] + inp[66] * layer_1_weights[19][66] + inp[67] * layer_1_weights[19][67] + inp[68] * layer_1_weights[19][68] + inp[69] * layer_1_weights[19][69] + inp[70] * layer_1_weights[19][70] + inp[71] * layer_1_weights[19][71] + inp[72] * layer_1_weights[19][72] + inp[73] * layer_1_weights[19][73] + inp[74] * layer_1_weights[19][74] + inp[75] * layer_1_weights[19][75] + inp[76] * layer_1_weights[19][76] + inp[77] * layer_1_weights[19][77] + inp[78] * layer_1_weights[19][78] + inp[79] * layer_1_weights[19][79] + inp[80] * layer_1_weights[19][80] + inp[81] * layer_1_weights[19][81] + inp[82] * layer_1_weights[19][82] + inp[83] * layer_1_weights[19][83] + inp[84] * layer_1_weights[19][84] + inp[85] * layer_1_weights[19][85] + inp[86] * layer_1_weights[19][86] + inp[87] * layer_1_weights[19][87] + inp[88] * layer_1_weights[19][88] + inp[89] * layer_1_weights[19][89] + inp[90] * layer_1_weights[19][90] + inp[91] * layer_1_weights[19][91] + inp[92] * layer_1_weights[19][92] + inp[93] * layer_1_weights[19][93] + inp[94] * layer_1_weights[19][94] + inp[95] * layer_1_weights[19][95] + inp[96] * layer_1_weights[19][96] + inp[97] * layer_1_weights[19][97] + inp[98] * layer_1_weights[19][98] + inp[99] * layer_1_weights[19][99] + inp[100] * layer_1_weights[19][100] + inp[101] * layer_1_weights[19][101] + inp[102] * layer_1_weights[19][102] + inp[103] * layer_1_weights[19][103] + inp[104] * layer_1_weights[19][104] + inp[105] * layer_1_weights[19][105] + inp[106] * layer_1_weights[19][106] + inp[107] * layer_1_weights[19][107] + inp[108] * layer_1_weights[19][108] + inp[109] * layer_1_weights[19][109] + inp[110] * layer_1_weights[19][110] + inp[111] * layer_1_weights[19][111] + inp[112] * layer_1_weights[19][112] + inp[113] * layer_1_weights[19][113] + inp[114] * layer_1_weights[19][114] + inp[115] * layer_1_weights[19][115] + inp[116] * layer_1_weights[19][116] + inp[117] * layer_1_weights[19][117] + inp[118] * layer_1_weights[19][118] + inp[119] * layer_1_weights[19][119] + inp[120] * layer_1_weights[19][120] + inp[121] * layer_1_weights[19][121] + inp[122] * layer_1_weights[19][122] + inp[123] * layer_1_weights[19][123] + inp[124] * layer_1_weights[19][124] + inp[125] * layer_1_weights[19][125] + inp[126] * layer_1_weights[19][126] + inp[127] * layer_1_weights[19][127] + inp[128] * layer_1_weights[19][128] + inp[129] * layer_1_weights[19][129] + inp[130] * layer_1_weights[19][130] + inp[131] * layer_1_weights[19][131] + inp[132] * layer_1_weights[19][132] + inp[133] * layer_1_weights[19][133] + inp[134] * layer_1_weights[19][134] + inp[135] * layer_1_weights[19][135] + inp[136] * layer_1_weights[19][136] + inp[137] * layer_1_weights[19][137] + inp[138] * layer_1_weights[19][138] + inp[139] * layer_1_weights[19][139] + inp[140] * layer_1_weights[19][140] + inp[141] * layer_1_weights[19][141] + inp[142] * layer_1_weights[19][142] + inp[143] * layer_1_weights[19][143]);
    assign layer_1_output_20 = relu(layer_1_biases[20] + inp[0] * layer_1_weights[20][0] + inp[1] * layer_1_weights[20][1] + inp[2] * layer_1_weights[20][2] + inp[3] * layer_1_weights[20][3] + inp[4] * layer_1_weights[20][4] + inp[5] * layer_1_weights[20][5] + inp[6] * layer_1_weights[20][6] + inp[7] * layer_1_weights[20][7] + inp[8] * layer_1_weights[20][8] + inp[9] * layer_1_weights[20][9] + inp[10] * layer_1_weights[20][10] + inp[11] * layer_1_weights[20][11] + inp[12] * layer_1_weights[20][12] + inp[13] * layer_1_weights[20][13] + inp[14] * layer_1_weights[20][14] + inp[15] * layer_1_weights[20][15] + inp[16] * layer_1_weights[20][16] + inp[17] * layer_1_weights[20][17] + inp[18] * layer_1_weights[20][18] + inp[19] * layer_1_weights[20][19] + inp[20] * layer_1_weights[20][20] + inp[21] * layer_1_weights[20][21] + inp[22] * layer_1_weights[20][22] + inp[23] * layer_1_weights[20][23] + inp[24] * layer_1_weights[20][24] + inp[25] * layer_1_weights[20][25] + inp[26] * layer_1_weights[20][26] + inp[27] * layer_1_weights[20][27] + inp[28] * layer_1_weights[20][28] + inp[29] * layer_1_weights[20][29] + inp[30] * layer_1_weights[20][30] + inp[31] * layer_1_weights[20][31] + inp[32] * layer_1_weights[20][32] + inp[33] * layer_1_weights[20][33] + inp[34] * layer_1_weights[20][34] + inp[35] * layer_1_weights[20][35] + inp[36] * layer_1_weights[20][36] + inp[37] * layer_1_weights[20][37] + inp[38] * layer_1_weights[20][38] + inp[39] * layer_1_weights[20][39] + inp[40] * layer_1_weights[20][40] + inp[41] * layer_1_weights[20][41] + inp[42] * layer_1_weights[20][42] + inp[43] * layer_1_weights[20][43] + inp[44] * layer_1_weights[20][44] + inp[45] * layer_1_weights[20][45] + inp[46] * layer_1_weights[20][46] + inp[47] * layer_1_weights[20][47] + inp[48] * layer_1_weights[20][48] + inp[49] * layer_1_weights[20][49] + inp[50] * layer_1_weights[20][50] + inp[51] * layer_1_weights[20][51] + inp[52] * layer_1_weights[20][52] + inp[53] * layer_1_weights[20][53] + inp[54] * layer_1_weights[20][54] + inp[55] * layer_1_weights[20][55] + inp[56] * layer_1_weights[20][56] + inp[57] * layer_1_weights[20][57] + inp[58] * layer_1_weights[20][58] + inp[59] * layer_1_weights[20][59] + inp[60] * layer_1_weights[20][60] + inp[61] * layer_1_weights[20][61] + inp[62] * layer_1_weights[20][62] + inp[63] * layer_1_weights[20][63] + inp[64] * layer_1_weights[20][64] + inp[65] * layer_1_weights[20][65] + inp[66] * layer_1_weights[20][66] + inp[67] * layer_1_weights[20][67] + inp[68] * layer_1_weights[20][68] + inp[69] * layer_1_weights[20][69] + inp[70] * layer_1_weights[20][70] + inp[71] * layer_1_weights[20][71] + inp[72] * layer_1_weights[20][72] + inp[73] * layer_1_weights[20][73] + inp[74] * layer_1_weights[20][74] + inp[75] * layer_1_weights[20][75] + inp[76] * layer_1_weights[20][76] + inp[77] * layer_1_weights[20][77] + inp[78] * layer_1_weights[20][78] + inp[79] * layer_1_weights[20][79] + inp[80] * layer_1_weights[20][80] + inp[81] * layer_1_weights[20][81] + inp[82] * layer_1_weights[20][82] + inp[83] * layer_1_weights[20][83] + inp[84] * layer_1_weights[20][84] + inp[85] * layer_1_weights[20][85] + inp[86] * layer_1_weights[20][86] + inp[87] * layer_1_weights[20][87] + inp[88] * layer_1_weights[20][88] + inp[89] * layer_1_weights[20][89] + inp[90] * layer_1_weights[20][90] + inp[91] * layer_1_weights[20][91] + inp[92] * layer_1_weights[20][92] + inp[93] * layer_1_weights[20][93] + inp[94] * layer_1_weights[20][94] + inp[95] * layer_1_weights[20][95] + inp[96] * layer_1_weights[20][96] + inp[97] * layer_1_weights[20][97] + inp[98] * layer_1_weights[20][98] + inp[99] * layer_1_weights[20][99] + inp[100] * layer_1_weights[20][100] + inp[101] * layer_1_weights[20][101] + inp[102] * layer_1_weights[20][102] + inp[103] * layer_1_weights[20][103] + inp[104] * layer_1_weights[20][104] + inp[105] * layer_1_weights[20][105] + inp[106] * layer_1_weights[20][106] + inp[107] * layer_1_weights[20][107] + inp[108] * layer_1_weights[20][108] + inp[109] * layer_1_weights[20][109] + inp[110] * layer_1_weights[20][110] + inp[111] * layer_1_weights[20][111] + inp[112] * layer_1_weights[20][112] + inp[113] * layer_1_weights[20][113] + inp[114] * layer_1_weights[20][114] + inp[115] * layer_1_weights[20][115] + inp[116] * layer_1_weights[20][116] + inp[117] * layer_1_weights[20][117] + inp[118] * layer_1_weights[20][118] + inp[119] * layer_1_weights[20][119] + inp[120] * layer_1_weights[20][120] + inp[121] * layer_1_weights[20][121] + inp[122] * layer_1_weights[20][122] + inp[123] * layer_1_weights[20][123] + inp[124] * layer_1_weights[20][124] + inp[125] * layer_1_weights[20][125] + inp[126] * layer_1_weights[20][126] + inp[127] * layer_1_weights[20][127] + inp[128] * layer_1_weights[20][128] + inp[129] * layer_1_weights[20][129] + inp[130] * layer_1_weights[20][130] + inp[131] * layer_1_weights[20][131] + inp[132] * layer_1_weights[20][132] + inp[133] * layer_1_weights[20][133] + inp[134] * layer_1_weights[20][134] + inp[135] * layer_1_weights[20][135] + inp[136] * layer_1_weights[20][136] + inp[137] * layer_1_weights[20][137] + inp[138] * layer_1_weights[20][138] + inp[139] * layer_1_weights[20][139] + inp[140] * layer_1_weights[20][140] + inp[141] * layer_1_weights[20][141] + inp[142] * layer_1_weights[20][142] + inp[143] * layer_1_weights[20][143]);
    assign layer_1_output_21 = relu(layer_1_biases[21] + inp[0] * layer_1_weights[21][0] + inp[1] * layer_1_weights[21][1] + inp[2] * layer_1_weights[21][2] + inp[3] * layer_1_weights[21][3] + inp[4] * layer_1_weights[21][4] + inp[5] * layer_1_weights[21][5] + inp[6] * layer_1_weights[21][6] + inp[7] * layer_1_weights[21][7] + inp[8] * layer_1_weights[21][8] + inp[9] * layer_1_weights[21][9] + inp[10] * layer_1_weights[21][10] + inp[11] * layer_1_weights[21][11] + inp[12] * layer_1_weights[21][12] + inp[13] * layer_1_weights[21][13] + inp[14] * layer_1_weights[21][14] + inp[15] * layer_1_weights[21][15] + inp[16] * layer_1_weights[21][16] + inp[17] * layer_1_weights[21][17] + inp[18] * layer_1_weights[21][18] + inp[19] * layer_1_weights[21][19] + inp[20] * layer_1_weights[21][20] + inp[21] * layer_1_weights[21][21] + inp[22] * layer_1_weights[21][22] + inp[23] * layer_1_weights[21][23] + inp[24] * layer_1_weights[21][24] + inp[25] * layer_1_weights[21][25] + inp[26] * layer_1_weights[21][26] + inp[27] * layer_1_weights[21][27] + inp[28] * layer_1_weights[21][28] + inp[29] * layer_1_weights[21][29] + inp[30] * layer_1_weights[21][30] + inp[31] * layer_1_weights[21][31] + inp[32] * layer_1_weights[21][32] + inp[33] * layer_1_weights[21][33] + inp[34] * layer_1_weights[21][34] + inp[35] * layer_1_weights[21][35] + inp[36] * layer_1_weights[21][36] + inp[37] * layer_1_weights[21][37] + inp[38] * layer_1_weights[21][38] + inp[39] * layer_1_weights[21][39] + inp[40] * layer_1_weights[21][40] + inp[41] * layer_1_weights[21][41] + inp[42] * layer_1_weights[21][42] + inp[43] * layer_1_weights[21][43] + inp[44] * layer_1_weights[21][44] + inp[45] * layer_1_weights[21][45] + inp[46] * layer_1_weights[21][46] + inp[47] * layer_1_weights[21][47] + inp[48] * layer_1_weights[21][48] + inp[49] * layer_1_weights[21][49] + inp[50] * layer_1_weights[21][50] + inp[51] * layer_1_weights[21][51] + inp[52] * layer_1_weights[21][52] + inp[53] * layer_1_weights[21][53] + inp[54] * layer_1_weights[21][54] + inp[55] * layer_1_weights[21][55] + inp[56] * layer_1_weights[21][56] + inp[57] * layer_1_weights[21][57] + inp[58] * layer_1_weights[21][58] + inp[59] * layer_1_weights[21][59] + inp[60] * layer_1_weights[21][60] + inp[61] * layer_1_weights[21][61] + inp[62] * layer_1_weights[21][62] + inp[63] * layer_1_weights[21][63] + inp[64] * layer_1_weights[21][64] + inp[65] * layer_1_weights[21][65] + inp[66] * layer_1_weights[21][66] + inp[67] * layer_1_weights[21][67] + inp[68] * layer_1_weights[21][68] + inp[69] * layer_1_weights[21][69] + inp[70] * layer_1_weights[21][70] + inp[71] * layer_1_weights[21][71] + inp[72] * layer_1_weights[21][72] + inp[73] * layer_1_weights[21][73] + inp[74] * layer_1_weights[21][74] + inp[75] * layer_1_weights[21][75] + inp[76] * layer_1_weights[21][76] + inp[77] * layer_1_weights[21][77] + inp[78] * layer_1_weights[21][78] + inp[79] * layer_1_weights[21][79] + inp[80] * layer_1_weights[21][80] + inp[81] * layer_1_weights[21][81] + inp[82] * layer_1_weights[21][82] + inp[83] * layer_1_weights[21][83] + inp[84] * layer_1_weights[21][84] + inp[85] * layer_1_weights[21][85] + inp[86] * layer_1_weights[21][86] + inp[87] * layer_1_weights[21][87] + inp[88] * layer_1_weights[21][88] + inp[89] * layer_1_weights[21][89] + inp[90] * layer_1_weights[21][90] + inp[91] * layer_1_weights[21][91] + inp[92] * layer_1_weights[21][92] + inp[93] * layer_1_weights[21][93] + inp[94] * layer_1_weights[21][94] + inp[95] * layer_1_weights[21][95] + inp[96] * layer_1_weights[21][96] + inp[97] * layer_1_weights[21][97] + inp[98] * layer_1_weights[21][98] + inp[99] * layer_1_weights[21][99] + inp[100] * layer_1_weights[21][100] + inp[101] * layer_1_weights[21][101] + inp[102] * layer_1_weights[21][102] + inp[103] * layer_1_weights[21][103] + inp[104] * layer_1_weights[21][104] + inp[105] * layer_1_weights[21][105] + inp[106] * layer_1_weights[21][106] + inp[107] * layer_1_weights[21][107] + inp[108] * layer_1_weights[21][108] + inp[109] * layer_1_weights[21][109] + inp[110] * layer_1_weights[21][110] + inp[111] * layer_1_weights[21][111] + inp[112] * layer_1_weights[21][112] + inp[113] * layer_1_weights[21][113] + inp[114] * layer_1_weights[21][114] + inp[115] * layer_1_weights[21][115] + inp[116] * layer_1_weights[21][116] + inp[117] * layer_1_weights[21][117] + inp[118] * layer_1_weights[21][118] + inp[119] * layer_1_weights[21][119] + inp[120] * layer_1_weights[21][120] + inp[121] * layer_1_weights[21][121] + inp[122] * layer_1_weights[21][122] + inp[123] * layer_1_weights[21][123] + inp[124] * layer_1_weights[21][124] + inp[125] * layer_1_weights[21][125] + inp[126] * layer_1_weights[21][126] + inp[127] * layer_1_weights[21][127] + inp[128] * layer_1_weights[21][128] + inp[129] * layer_1_weights[21][129] + inp[130] * layer_1_weights[21][130] + inp[131] * layer_1_weights[21][131] + inp[132] * layer_1_weights[21][132] + inp[133] * layer_1_weights[21][133] + inp[134] * layer_1_weights[21][134] + inp[135] * layer_1_weights[21][135] + inp[136] * layer_1_weights[21][136] + inp[137] * layer_1_weights[21][137] + inp[138] * layer_1_weights[21][138] + inp[139] * layer_1_weights[21][139] + inp[140] * layer_1_weights[21][140] + inp[141] * layer_1_weights[21][141] + inp[142] * layer_1_weights[21][142] + inp[143] * layer_1_weights[21][143]);
    assign layer_1_output_22 = relu(layer_1_biases[22] + inp[0] * layer_1_weights[22][0] + inp[1] * layer_1_weights[22][1] + inp[2] * layer_1_weights[22][2] + inp[3] * layer_1_weights[22][3] + inp[4] * layer_1_weights[22][4] + inp[5] * layer_1_weights[22][5] + inp[6] * layer_1_weights[22][6] + inp[7] * layer_1_weights[22][7] + inp[8] * layer_1_weights[22][8] + inp[9] * layer_1_weights[22][9] + inp[10] * layer_1_weights[22][10] + inp[11] * layer_1_weights[22][11] + inp[12] * layer_1_weights[22][12] + inp[13] * layer_1_weights[22][13] + inp[14] * layer_1_weights[22][14] + inp[15] * layer_1_weights[22][15] + inp[16] * layer_1_weights[22][16] + inp[17] * layer_1_weights[22][17] + inp[18] * layer_1_weights[22][18] + inp[19] * layer_1_weights[22][19] + inp[20] * layer_1_weights[22][20] + inp[21] * layer_1_weights[22][21] + inp[22] * layer_1_weights[22][22] + inp[23] * layer_1_weights[22][23] + inp[24] * layer_1_weights[22][24] + inp[25] * layer_1_weights[22][25] + inp[26] * layer_1_weights[22][26] + inp[27] * layer_1_weights[22][27] + inp[28] * layer_1_weights[22][28] + inp[29] * layer_1_weights[22][29] + inp[30] * layer_1_weights[22][30] + inp[31] * layer_1_weights[22][31] + inp[32] * layer_1_weights[22][32] + inp[33] * layer_1_weights[22][33] + inp[34] * layer_1_weights[22][34] + inp[35] * layer_1_weights[22][35] + inp[36] * layer_1_weights[22][36] + inp[37] * layer_1_weights[22][37] + inp[38] * layer_1_weights[22][38] + inp[39] * layer_1_weights[22][39] + inp[40] * layer_1_weights[22][40] + inp[41] * layer_1_weights[22][41] + inp[42] * layer_1_weights[22][42] + inp[43] * layer_1_weights[22][43] + inp[44] * layer_1_weights[22][44] + inp[45] * layer_1_weights[22][45] + inp[46] * layer_1_weights[22][46] + inp[47] * layer_1_weights[22][47] + inp[48] * layer_1_weights[22][48] + inp[49] * layer_1_weights[22][49] + inp[50] * layer_1_weights[22][50] + inp[51] * layer_1_weights[22][51] + inp[52] * layer_1_weights[22][52] + inp[53] * layer_1_weights[22][53] + inp[54] * layer_1_weights[22][54] + inp[55] * layer_1_weights[22][55] + inp[56] * layer_1_weights[22][56] + inp[57] * layer_1_weights[22][57] + inp[58] * layer_1_weights[22][58] + inp[59] * layer_1_weights[22][59] + inp[60] * layer_1_weights[22][60] + inp[61] * layer_1_weights[22][61] + inp[62] * layer_1_weights[22][62] + inp[63] * layer_1_weights[22][63] + inp[64] * layer_1_weights[22][64] + inp[65] * layer_1_weights[22][65] + inp[66] * layer_1_weights[22][66] + inp[67] * layer_1_weights[22][67] + inp[68] * layer_1_weights[22][68] + inp[69] * layer_1_weights[22][69] + inp[70] * layer_1_weights[22][70] + inp[71] * layer_1_weights[22][71] + inp[72] * layer_1_weights[22][72] + inp[73] * layer_1_weights[22][73] + inp[74] * layer_1_weights[22][74] + inp[75] * layer_1_weights[22][75] + inp[76] * layer_1_weights[22][76] + inp[77] * layer_1_weights[22][77] + inp[78] * layer_1_weights[22][78] + inp[79] * layer_1_weights[22][79] + inp[80] * layer_1_weights[22][80] + inp[81] * layer_1_weights[22][81] + inp[82] * layer_1_weights[22][82] + inp[83] * layer_1_weights[22][83] + inp[84] * layer_1_weights[22][84] + inp[85] * layer_1_weights[22][85] + inp[86] * layer_1_weights[22][86] + inp[87] * layer_1_weights[22][87] + inp[88] * layer_1_weights[22][88] + inp[89] * layer_1_weights[22][89] + inp[90] * layer_1_weights[22][90] + inp[91] * layer_1_weights[22][91] + inp[92] * layer_1_weights[22][92] + inp[93] * layer_1_weights[22][93] + inp[94] * layer_1_weights[22][94] + inp[95] * layer_1_weights[22][95] + inp[96] * layer_1_weights[22][96] + inp[97] * layer_1_weights[22][97] + inp[98] * layer_1_weights[22][98] + inp[99] * layer_1_weights[22][99] + inp[100] * layer_1_weights[22][100] + inp[101] * layer_1_weights[22][101] + inp[102] * layer_1_weights[22][102] + inp[103] * layer_1_weights[22][103] + inp[104] * layer_1_weights[22][104] + inp[105] * layer_1_weights[22][105] + inp[106] * layer_1_weights[22][106] + inp[107] * layer_1_weights[22][107] + inp[108] * layer_1_weights[22][108] + inp[109] * layer_1_weights[22][109] + inp[110] * layer_1_weights[22][110] + inp[111] * layer_1_weights[22][111] + inp[112] * layer_1_weights[22][112] + inp[113] * layer_1_weights[22][113] + inp[114] * layer_1_weights[22][114] + inp[115] * layer_1_weights[22][115] + inp[116] * layer_1_weights[22][116] + inp[117] * layer_1_weights[22][117] + inp[118] * layer_1_weights[22][118] + inp[119] * layer_1_weights[22][119] + inp[120] * layer_1_weights[22][120] + inp[121] * layer_1_weights[22][121] + inp[122] * layer_1_weights[22][122] + inp[123] * layer_1_weights[22][123] + inp[124] * layer_1_weights[22][124] + inp[125] * layer_1_weights[22][125] + inp[126] * layer_1_weights[22][126] + inp[127] * layer_1_weights[22][127] + inp[128] * layer_1_weights[22][128] + inp[129] * layer_1_weights[22][129] + inp[130] * layer_1_weights[22][130] + inp[131] * layer_1_weights[22][131] + inp[132] * layer_1_weights[22][132] + inp[133] * layer_1_weights[22][133] + inp[134] * layer_1_weights[22][134] + inp[135] * layer_1_weights[22][135] + inp[136] * layer_1_weights[22][136] + inp[137] * layer_1_weights[22][137] + inp[138] * layer_1_weights[22][138] + inp[139] * layer_1_weights[22][139] + inp[140] * layer_1_weights[22][140] + inp[141] * layer_1_weights[22][141] + inp[142] * layer_1_weights[22][142] + inp[143] * layer_1_weights[22][143]);
    assign layer_1_output_23 = relu(layer_1_biases[23] + inp[0] * layer_1_weights[23][0] + inp[1] * layer_1_weights[23][1] + inp[2] * layer_1_weights[23][2] + inp[3] * layer_1_weights[23][3] + inp[4] * layer_1_weights[23][4] + inp[5] * layer_1_weights[23][5] + inp[6] * layer_1_weights[23][6] + inp[7] * layer_1_weights[23][7] + inp[8] * layer_1_weights[23][8] + inp[9] * layer_1_weights[23][9] + inp[10] * layer_1_weights[23][10] + inp[11] * layer_1_weights[23][11] + inp[12] * layer_1_weights[23][12] + inp[13] * layer_1_weights[23][13] + inp[14] * layer_1_weights[23][14] + inp[15] * layer_1_weights[23][15] + inp[16] * layer_1_weights[23][16] + inp[17] * layer_1_weights[23][17] + inp[18] * layer_1_weights[23][18] + inp[19] * layer_1_weights[23][19] + inp[20] * layer_1_weights[23][20] + inp[21] * layer_1_weights[23][21] + inp[22] * layer_1_weights[23][22] + inp[23] * layer_1_weights[23][23] + inp[24] * layer_1_weights[23][24] + inp[25] * layer_1_weights[23][25] + inp[26] * layer_1_weights[23][26] + inp[27] * layer_1_weights[23][27] + inp[28] * layer_1_weights[23][28] + inp[29] * layer_1_weights[23][29] + inp[30] * layer_1_weights[23][30] + inp[31] * layer_1_weights[23][31] + inp[32] * layer_1_weights[23][32] + inp[33] * layer_1_weights[23][33] + inp[34] * layer_1_weights[23][34] + inp[35] * layer_1_weights[23][35] + inp[36] * layer_1_weights[23][36] + inp[37] * layer_1_weights[23][37] + inp[38] * layer_1_weights[23][38] + inp[39] * layer_1_weights[23][39] + inp[40] * layer_1_weights[23][40] + inp[41] * layer_1_weights[23][41] + inp[42] * layer_1_weights[23][42] + inp[43] * layer_1_weights[23][43] + inp[44] * layer_1_weights[23][44] + inp[45] * layer_1_weights[23][45] + inp[46] * layer_1_weights[23][46] + inp[47] * layer_1_weights[23][47] + inp[48] * layer_1_weights[23][48] + inp[49] * layer_1_weights[23][49] + inp[50] * layer_1_weights[23][50] + inp[51] * layer_1_weights[23][51] + inp[52] * layer_1_weights[23][52] + inp[53] * layer_1_weights[23][53] + inp[54] * layer_1_weights[23][54] + inp[55] * layer_1_weights[23][55] + inp[56] * layer_1_weights[23][56] + inp[57] * layer_1_weights[23][57] + inp[58] * layer_1_weights[23][58] + inp[59] * layer_1_weights[23][59] + inp[60] * layer_1_weights[23][60] + inp[61] * layer_1_weights[23][61] + inp[62] * layer_1_weights[23][62] + inp[63] * layer_1_weights[23][63] + inp[64] * layer_1_weights[23][64] + inp[65] * layer_1_weights[23][65] + inp[66] * layer_1_weights[23][66] + inp[67] * layer_1_weights[23][67] + inp[68] * layer_1_weights[23][68] + inp[69] * layer_1_weights[23][69] + inp[70] * layer_1_weights[23][70] + inp[71] * layer_1_weights[23][71] + inp[72] * layer_1_weights[23][72] + inp[73] * layer_1_weights[23][73] + inp[74] * layer_1_weights[23][74] + inp[75] * layer_1_weights[23][75] + inp[76] * layer_1_weights[23][76] + inp[77] * layer_1_weights[23][77] + inp[78] * layer_1_weights[23][78] + inp[79] * layer_1_weights[23][79] + inp[80] * layer_1_weights[23][80] + inp[81] * layer_1_weights[23][81] + inp[82] * layer_1_weights[23][82] + inp[83] * layer_1_weights[23][83] + inp[84] * layer_1_weights[23][84] + inp[85] * layer_1_weights[23][85] + inp[86] * layer_1_weights[23][86] + inp[87] * layer_1_weights[23][87] + inp[88] * layer_1_weights[23][88] + inp[89] * layer_1_weights[23][89] + inp[90] * layer_1_weights[23][90] + inp[91] * layer_1_weights[23][91] + inp[92] * layer_1_weights[23][92] + inp[93] * layer_1_weights[23][93] + inp[94] * layer_1_weights[23][94] + inp[95] * layer_1_weights[23][95] + inp[96] * layer_1_weights[23][96] + inp[97] * layer_1_weights[23][97] + inp[98] * layer_1_weights[23][98] + inp[99] * layer_1_weights[23][99] + inp[100] * layer_1_weights[23][100] + inp[101] * layer_1_weights[23][101] + inp[102] * layer_1_weights[23][102] + inp[103] * layer_1_weights[23][103] + inp[104] * layer_1_weights[23][104] + inp[105] * layer_1_weights[23][105] + inp[106] * layer_1_weights[23][106] + inp[107] * layer_1_weights[23][107] + inp[108] * layer_1_weights[23][108] + inp[109] * layer_1_weights[23][109] + inp[110] * layer_1_weights[23][110] + inp[111] * layer_1_weights[23][111] + inp[112] * layer_1_weights[23][112] + inp[113] * layer_1_weights[23][113] + inp[114] * layer_1_weights[23][114] + inp[115] * layer_1_weights[23][115] + inp[116] * layer_1_weights[23][116] + inp[117] * layer_1_weights[23][117] + inp[118] * layer_1_weights[23][118] + inp[119] * layer_1_weights[23][119] + inp[120] * layer_1_weights[23][120] + inp[121] * layer_1_weights[23][121] + inp[122] * layer_1_weights[23][122] + inp[123] * layer_1_weights[23][123] + inp[124] * layer_1_weights[23][124] + inp[125] * layer_1_weights[23][125] + inp[126] * layer_1_weights[23][126] + inp[127] * layer_1_weights[23][127] + inp[128] * layer_1_weights[23][128] + inp[129] * layer_1_weights[23][129] + inp[130] * layer_1_weights[23][130] + inp[131] * layer_1_weights[23][131] + inp[132] * layer_1_weights[23][132] + inp[133] * layer_1_weights[23][133] + inp[134] * layer_1_weights[23][134] + inp[135] * layer_1_weights[23][135] + inp[136] * layer_1_weights[23][136] + inp[137] * layer_1_weights[23][137] + inp[138] * layer_1_weights[23][138] + inp[139] * layer_1_weights[23][139] + inp[140] * layer_1_weights[23][140] + inp[141] * layer_1_weights[23][141] + inp[142] * layer_1_weights[23][142] + inp[143] * layer_1_weights[23][143]);
    assign layer_1_output_24 = relu(layer_1_biases[24] + inp[0] * layer_1_weights[24][0] + inp[1] * layer_1_weights[24][1] + inp[2] * layer_1_weights[24][2] + inp[3] * layer_1_weights[24][3] + inp[4] * layer_1_weights[24][4] + inp[5] * layer_1_weights[24][5] + inp[6] * layer_1_weights[24][6] + inp[7] * layer_1_weights[24][7] + inp[8] * layer_1_weights[24][8] + inp[9] * layer_1_weights[24][9] + inp[10] * layer_1_weights[24][10] + inp[11] * layer_1_weights[24][11] + inp[12] * layer_1_weights[24][12] + inp[13] * layer_1_weights[24][13] + inp[14] * layer_1_weights[24][14] + inp[15] * layer_1_weights[24][15] + inp[16] * layer_1_weights[24][16] + inp[17] * layer_1_weights[24][17] + inp[18] * layer_1_weights[24][18] + inp[19] * layer_1_weights[24][19] + inp[20] * layer_1_weights[24][20] + inp[21] * layer_1_weights[24][21] + inp[22] * layer_1_weights[24][22] + inp[23] * layer_1_weights[24][23] + inp[24] * layer_1_weights[24][24] + inp[25] * layer_1_weights[24][25] + inp[26] * layer_1_weights[24][26] + inp[27] * layer_1_weights[24][27] + inp[28] * layer_1_weights[24][28] + inp[29] * layer_1_weights[24][29] + inp[30] * layer_1_weights[24][30] + inp[31] * layer_1_weights[24][31] + inp[32] * layer_1_weights[24][32] + inp[33] * layer_1_weights[24][33] + inp[34] * layer_1_weights[24][34] + inp[35] * layer_1_weights[24][35] + inp[36] * layer_1_weights[24][36] + inp[37] * layer_1_weights[24][37] + inp[38] * layer_1_weights[24][38] + inp[39] * layer_1_weights[24][39] + inp[40] * layer_1_weights[24][40] + inp[41] * layer_1_weights[24][41] + inp[42] * layer_1_weights[24][42] + inp[43] * layer_1_weights[24][43] + inp[44] * layer_1_weights[24][44] + inp[45] * layer_1_weights[24][45] + inp[46] * layer_1_weights[24][46] + inp[47] * layer_1_weights[24][47] + inp[48] * layer_1_weights[24][48] + inp[49] * layer_1_weights[24][49] + inp[50] * layer_1_weights[24][50] + inp[51] * layer_1_weights[24][51] + inp[52] * layer_1_weights[24][52] + inp[53] * layer_1_weights[24][53] + inp[54] * layer_1_weights[24][54] + inp[55] * layer_1_weights[24][55] + inp[56] * layer_1_weights[24][56] + inp[57] * layer_1_weights[24][57] + inp[58] * layer_1_weights[24][58] + inp[59] * layer_1_weights[24][59] + inp[60] * layer_1_weights[24][60] + inp[61] * layer_1_weights[24][61] + inp[62] * layer_1_weights[24][62] + inp[63] * layer_1_weights[24][63] + inp[64] * layer_1_weights[24][64] + inp[65] * layer_1_weights[24][65] + inp[66] * layer_1_weights[24][66] + inp[67] * layer_1_weights[24][67] + inp[68] * layer_1_weights[24][68] + inp[69] * layer_1_weights[24][69] + inp[70] * layer_1_weights[24][70] + inp[71] * layer_1_weights[24][71] + inp[72] * layer_1_weights[24][72] + inp[73] * layer_1_weights[24][73] + inp[74] * layer_1_weights[24][74] + inp[75] * layer_1_weights[24][75] + inp[76] * layer_1_weights[24][76] + inp[77] * layer_1_weights[24][77] + inp[78] * layer_1_weights[24][78] + inp[79] * layer_1_weights[24][79] + inp[80] * layer_1_weights[24][80] + inp[81] * layer_1_weights[24][81] + inp[82] * layer_1_weights[24][82] + inp[83] * layer_1_weights[24][83] + inp[84] * layer_1_weights[24][84] + inp[85] * layer_1_weights[24][85] + inp[86] * layer_1_weights[24][86] + inp[87] * layer_1_weights[24][87] + inp[88] * layer_1_weights[24][88] + inp[89] * layer_1_weights[24][89] + inp[90] * layer_1_weights[24][90] + inp[91] * layer_1_weights[24][91] + inp[92] * layer_1_weights[24][92] + inp[93] * layer_1_weights[24][93] + inp[94] * layer_1_weights[24][94] + inp[95] * layer_1_weights[24][95] + inp[96] * layer_1_weights[24][96] + inp[97] * layer_1_weights[24][97] + inp[98] * layer_1_weights[24][98] + inp[99] * layer_1_weights[24][99] + inp[100] * layer_1_weights[24][100] + inp[101] * layer_1_weights[24][101] + inp[102] * layer_1_weights[24][102] + inp[103] * layer_1_weights[24][103] + inp[104] * layer_1_weights[24][104] + inp[105] * layer_1_weights[24][105] + inp[106] * layer_1_weights[24][106] + inp[107] * layer_1_weights[24][107] + inp[108] * layer_1_weights[24][108] + inp[109] * layer_1_weights[24][109] + inp[110] * layer_1_weights[24][110] + inp[111] * layer_1_weights[24][111] + inp[112] * layer_1_weights[24][112] + inp[113] * layer_1_weights[24][113] + inp[114] * layer_1_weights[24][114] + inp[115] * layer_1_weights[24][115] + inp[116] * layer_1_weights[24][116] + inp[117] * layer_1_weights[24][117] + inp[118] * layer_1_weights[24][118] + inp[119] * layer_1_weights[24][119] + inp[120] * layer_1_weights[24][120] + inp[121] * layer_1_weights[24][121] + inp[122] * layer_1_weights[24][122] + inp[123] * layer_1_weights[24][123] + inp[124] * layer_1_weights[24][124] + inp[125] * layer_1_weights[24][125] + inp[126] * layer_1_weights[24][126] + inp[127] * layer_1_weights[24][127] + inp[128] * layer_1_weights[24][128] + inp[129] * layer_1_weights[24][129] + inp[130] * layer_1_weights[24][130] + inp[131] * layer_1_weights[24][131] + inp[132] * layer_1_weights[24][132] + inp[133] * layer_1_weights[24][133] + inp[134] * layer_1_weights[24][134] + inp[135] * layer_1_weights[24][135] + inp[136] * layer_1_weights[24][136] + inp[137] * layer_1_weights[24][137] + inp[138] * layer_1_weights[24][138] + inp[139] * layer_1_weights[24][139] + inp[140] * layer_1_weights[24][140] + inp[141] * layer_1_weights[24][141] + inp[142] * layer_1_weights[24][142] + inp[143] * layer_1_weights[24][143]);
    assign layer_1_output_25 = relu(layer_1_biases[25] + inp[0] * layer_1_weights[25][0] + inp[1] * layer_1_weights[25][1] + inp[2] * layer_1_weights[25][2] + inp[3] * layer_1_weights[25][3] + inp[4] * layer_1_weights[25][4] + inp[5] * layer_1_weights[25][5] + inp[6] * layer_1_weights[25][6] + inp[7] * layer_1_weights[25][7] + inp[8] * layer_1_weights[25][8] + inp[9] * layer_1_weights[25][9] + inp[10] * layer_1_weights[25][10] + inp[11] * layer_1_weights[25][11] + inp[12] * layer_1_weights[25][12] + inp[13] * layer_1_weights[25][13] + inp[14] * layer_1_weights[25][14] + inp[15] * layer_1_weights[25][15] + inp[16] * layer_1_weights[25][16] + inp[17] * layer_1_weights[25][17] + inp[18] * layer_1_weights[25][18] + inp[19] * layer_1_weights[25][19] + inp[20] * layer_1_weights[25][20] + inp[21] * layer_1_weights[25][21] + inp[22] * layer_1_weights[25][22] + inp[23] * layer_1_weights[25][23] + inp[24] * layer_1_weights[25][24] + inp[25] * layer_1_weights[25][25] + inp[26] * layer_1_weights[25][26] + inp[27] * layer_1_weights[25][27] + inp[28] * layer_1_weights[25][28] + inp[29] * layer_1_weights[25][29] + inp[30] * layer_1_weights[25][30] + inp[31] * layer_1_weights[25][31] + inp[32] * layer_1_weights[25][32] + inp[33] * layer_1_weights[25][33] + inp[34] * layer_1_weights[25][34] + inp[35] * layer_1_weights[25][35] + inp[36] * layer_1_weights[25][36] + inp[37] * layer_1_weights[25][37] + inp[38] * layer_1_weights[25][38] + inp[39] * layer_1_weights[25][39] + inp[40] * layer_1_weights[25][40] + inp[41] * layer_1_weights[25][41] + inp[42] * layer_1_weights[25][42] + inp[43] * layer_1_weights[25][43] + inp[44] * layer_1_weights[25][44] + inp[45] * layer_1_weights[25][45] + inp[46] * layer_1_weights[25][46] + inp[47] * layer_1_weights[25][47] + inp[48] * layer_1_weights[25][48] + inp[49] * layer_1_weights[25][49] + inp[50] * layer_1_weights[25][50] + inp[51] * layer_1_weights[25][51] + inp[52] * layer_1_weights[25][52] + inp[53] * layer_1_weights[25][53] + inp[54] * layer_1_weights[25][54] + inp[55] * layer_1_weights[25][55] + inp[56] * layer_1_weights[25][56] + inp[57] * layer_1_weights[25][57] + inp[58] * layer_1_weights[25][58] + inp[59] * layer_1_weights[25][59] + inp[60] * layer_1_weights[25][60] + inp[61] * layer_1_weights[25][61] + inp[62] * layer_1_weights[25][62] + inp[63] * layer_1_weights[25][63] + inp[64] * layer_1_weights[25][64] + inp[65] * layer_1_weights[25][65] + inp[66] * layer_1_weights[25][66] + inp[67] * layer_1_weights[25][67] + inp[68] * layer_1_weights[25][68] + inp[69] * layer_1_weights[25][69] + inp[70] * layer_1_weights[25][70] + inp[71] * layer_1_weights[25][71] + inp[72] * layer_1_weights[25][72] + inp[73] * layer_1_weights[25][73] + inp[74] * layer_1_weights[25][74] + inp[75] * layer_1_weights[25][75] + inp[76] * layer_1_weights[25][76] + inp[77] * layer_1_weights[25][77] + inp[78] * layer_1_weights[25][78] + inp[79] * layer_1_weights[25][79] + inp[80] * layer_1_weights[25][80] + inp[81] * layer_1_weights[25][81] + inp[82] * layer_1_weights[25][82] + inp[83] * layer_1_weights[25][83] + inp[84] * layer_1_weights[25][84] + inp[85] * layer_1_weights[25][85] + inp[86] * layer_1_weights[25][86] + inp[87] * layer_1_weights[25][87] + inp[88] * layer_1_weights[25][88] + inp[89] * layer_1_weights[25][89] + inp[90] * layer_1_weights[25][90] + inp[91] * layer_1_weights[25][91] + inp[92] * layer_1_weights[25][92] + inp[93] * layer_1_weights[25][93] + inp[94] * layer_1_weights[25][94] + inp[95] * layer_1_weights[25][95] + inp[96] * layer_1_weights[25][96] + inp[97] * layer_1_weights[25][97] + inp[98] * layer_1_weights[25][98] + inp[99] * layer_1_weights[25][99] + inp[100] * layer_1_weights[25][100] + inp[101] * layer_1_weights[25][101] + inp[102] * layer_1_weights[25][102] + inp[103] * layer_1_weights[25][103] + inp[104] * layer_1_weights[25][104] + inp[105] * layer_1_weights[25][105] + inp[106] * layer_1_weights[25][106] + inp[107] * layer_1_weights[25][107] + inp[108] * layer_1_weights[25][108] + inp[109] * layer_1_weights[25][109] + inp[110] * layer_1_weights[25][110] + inp[111] * layer_1_weights[25][111] + inp[112] * layer_1_weights[25][112] + inp[113] * layer_1_weights[25][113] + inp[114] * layer_1_weights[25][114] + inp[115] * layer_1_weights[25][115] + inp[116] * layer_1_weights[25][116] + inp[117] * layer_1_weights[25][117] + inp[118] * layer_1_weights[25][118] + inp[119] * layer_1_weights[25][119] + inp[120] * layer_1_weights[25][120] + inp[121] * layer_1_weights[25][121] + inp[122] * layer_1_weights[25][122] + inp[123] * layer_1_weights[25][123] + inp[124] * layer_1_weights[25][124] + inp[125] * layer_1_weights[25][125] + inp[126] * layer_1_weights[25][126] + inp[127] * layer_1_weights[25][127] + inp[128] * layer_1_weights[25][128] + inp[129] * layer_1_weights[25][129] + inp[130] * layer_1_weights[25][130] + inp[131] * layer_1_weights[25][131] + inp[132] * layer_1_weights[25][132] + inp[133] * layer_1_weights[25][133] + inp[134] * layer_1_weights[25][134] + inp[135] * layer_1_weights[25][135] + inp[136] * layer_1_weights[25][136] + inp[137] * layer_1_weights[25][137] + inp[138] * layer_1_weights[25][138] + inp[139] * layer_1_weights[25][139] + inp[140] * layer_1_weights[25][140] + inp[141] * layer_1_weights[25][141] + inp[142] * layer_1_weights[25][142] + inp[143] * layer_1_weights[25][143]);
    assign layer_1_output_26 = relu(layer_1_biases[26] + inp[0] * layer_1_weights[26][0] + inp[1] * layer_1_weights[26][1] + inp[2] * layer_1_weights[26][2] + inp[3] * layer_1_weights[26][3] + inp[4] * layer_1_weights[26][4] + inp[5] * layer_1_weights[26][5] + inp[6] * layer_1_weights[26][6] + inp[7] * layer_1_weights[26][7] + inp[8] * layer_1_weights[26][8] + inp[9] * layer_1_weights[26][9] + inp[10] * layer_1_weights[26][10] + inp[11] * layer_1_weights[26][11] + inp[12] * layer_1_weights[26][12] + inp[13] * layer_1_weights[26][13] + inp[14] * layer_1_weights[26][14] + inp[15] * layer_1_weights[26][15] + inp[16] * layer_1_weights[26][16] + inp[17] * layer_1_weights[26][17] + inp[18] * layer_1_weights[26][18] + inp[19] * layer_1_weights[26][19] + inp[20] * layer_1_weights[26][20] + inp[21] * layer_1_weights[26][21] + inp[22] * layer_1_weights[26][22] + inp[23] * layer_1_weights[26][23] + inp[24] * layer_1_weights[26][24] + inp[25] * layer_1_weights[26][25] + inp[26] * layer_1_weights[26][26] + inp[27] * layer_1_weights[26][27] + inp[28] * layer_1_weights[26][28] + inp[29] * layer_1_weights[26][29] + inp[30] * layer_1_weights[26][30] + inp[31] * layer_1_weights[26][31] + inp[32] * layer_1_weights[26][32] + inp[33] * layer_1_weights[26][33] + inp[34] * layer_1_weights[26][34] + inp[35] * layer_1_weights[26][35] + inp[36] * layer_1_weights[26][36] + inp[37] * layer_1_weights[26][37] + inp[38] * layer_1_weights[26][38] + inp[39] * layer_1_weights[26][39] + inp[40] * layer_1_weights[26][40] + inp[41] * layer_1_weights[26][41] + inp[42] * layer_1_weights[26][42] + inp[43] * layer_1_weights[26][43] + inp[44] * layer_1_weights[26][44] + inp[45] * layer_1_weights[26][45] + inp[46] * layer_1_weights[26][46] + inp[47] * layer_1_weights[26][47] + inp[48] * layer_1_weights[26][48] + inp[49] * layer_1_weights[26][49] + inp[50] * layer_1_weights[26][50] + inp[51] * layer_1_weights[26][51] + inp[52] * layer_1_weights[26][52] + inp[53] * layer_1_weights[26][53] + inp[54] * layer_1_weights[26][54] + inp[55] * layer_1_weights[26][55] + inp[56] * layer_1_weights[26][56] + inp[57] * layer_1_weights[26][57] + inp[58] * layer_1_weights[26][58] + inp[59] * layer_1_weights[26][59] + inp[60] * layer_1_weights[26][60] + inp[61] * layer_1_weights[26][61] + inp[62] * layer_1_weights[26][62] + inp[63] * layer_1_weights[26][63] + inp[64] * layer_1_weights[26][64] + inp[65] * layer_1_weights[26][65] + inp[66] * layer_1_weights[26][66] + inp[67] * layer_1_weights[26][67] + inp[68] * layer_1_weights[26][68] + inp[69] * layer_1_weights[26][69] + inp[70] * layer_1_weights[26][70] + inp[71] * layer_1_weights[26][71] + inp[72] * layer_1_weights[26][72] + inp[73] * layer_1_weights[26][73] + inp[74] * layer_1_weights[26][74] + inp[75] * layer_1_weights[26][75] + inp[76] * layer_1_weights[26][76] + inp[77] * layer_1_weights[26][77] + inp[78] * layer_1_weights[26][78] + inp[79] * layer_1_weights[26][79] + inp[80] * layer_1_weights[26][80] + inp[81] * layer_1_weights[26][81] + inp[82] * layer_1_weights[26][82] + inp[83] * layer_1_weights[26][83] + inp[84] * layer_1_weights[26][84] + inp[85] * layer_1_weights[26][85] + inp[86] * layer_1_weights[26][86] + inp[87] * layer_1_weights[26][87] + inp[88] * layer_1_weights[26][88] + inp[89] * layer_1_weights[26][89] + inp[90] * layer_1_weights[26][90] + inp[91] * layer_1_weights[26][91] + inp[92] * layer_1_weights[26][92] + inp[93] * layer_1_weights[26][93] + inp[94] * layer_1_weights[26][94] + inp[95] * layer_1_weights[26][95] + inp[96] * layer_1_weights[26][96] + inp[97] * layer_1_weights[26][97] + inp[98] * layer_1_weights[26][98] + inp[99] * layer_1_weights[26][99] + inp[100] * layer_1_weights[26][100] + inp[101] * layer_1_weights[26][101] + inp[102] * layer_1_weights[26][102] + inp[103] * layer_1_weights[26][103] + inp[104] * layer_1_weights[26][104] + inp[105] * layer_1_weights[26][105] + inp[106] * layer_1_weights[26][106] + inp[107] * layer_1_weights[26][107] + inp[108] * layer_1_weights[26][108] + inp[109] * layer_1_weights[26][109] + inp[110] * layer_1_weights[26][110] + inp[111] * layer_1_weights[26][111] + inp[112] * layer_1_weights[26][112] + inp[113] * layer_1_weights[26][113] + inp[114] * layer_1_weights[26][114] + inp[115] * layer_1_weights[26][115] + inp[116] * layer_1_weights[26][116] + inp[117] * layer_1_weights[26][117] + inp[118] * layer_1_weights[26][118] + inp[119] * layer_1_weights[26][119] + inp[120] * layer_1_weights[26][120] + inp[121] * layer_1_weights[26][121] + inp[122] * layer_1_weights[26][122] + inp[123] * layer_1_weights[26][123] + inp[124] * layer_1_weights[26][124] + inp[125] * layer_1_weights[26][125] + inp[126] * layer_1_weights[26][126] + inp[127] * layer_1_weights[26][127] + inp[128] * layer_1_weights[26][128] + inp[129] * layer_1_weights[26][129] + inp[130] * layer_1_weights[26][130] + inp[131] * layer_1_weights[26][131] + inp[132] * layer_1_weights[26][132] + inp[133] * layer_1_weights[26][133] + inp[134] * layer_1_weights[26][134] + inp[135] * layer_1_weights[26][135] + inp[136] * layer_1_weights[26][136] + inp[137] * layer_1_weights[26][137] + inp[138] * layer_1_weights[26][138] + inp[139] * layer_1_weights[26][139] + inp[140] * layer_1_weights[26][140] + inp[141] * layer_1_weights[26][141] + inp[142] * layer_1_weights[26][142] + inp[143] * layer_1_weights[26][143]);
    assign layer_1_output_27 = relu(layer_1_biases[27] + inp[0] * layer_1_weights[27][0] + inp[1] * layer_1_weights[27][1] + inp[2] * layer_1_weights[27][2] + inp[3] * layer_1_weights[27][3] + inp[4] * layer_1_weights[27][4] + inp[5] * layer_1_weights[27][5] + inp[6] * layer_1_weights[27][6] + inp[7] * layer_1_weights[27][7] + inp[8] * layer_1_weights[27][8] + inp[9] * layer_1_weights[27][9] + inp[10] * layer_1_weights[27][10] + inp[11] * layer_1_weights[27][11] + inp[12] * layer_1_weights[27][12] + inp[13] * layer_1_weights[27][13] + inp[14] * layer_1_weights[27][14] + inp[15] * layer_1_weights[27][15] + inp[16] * layer_1_weights[27][16] + inp[17] * layer_1_weights[27][17] + inp[18] * layer_1_weights[27][18] + inp[19] * layer_1_weights[27][19] + inp[20] * layer_1_weights[27][20] + inp[21] * layer_1_weights[27][21] + inp[22] * layer_1_weights[27][22] + inp[23] * layer_1_weights[27][23] + inp[24] * layer_1_weights[27][24] + inp[25] * layer_1_weights[27][25] + inp[26] * layer_1_weights[27][26] + inp[27] * layer_1_weights[27][27] + inp[28] * layer_1_weights[27][28] + inp[29] * layer_1_weights[27][29] + inp[30] * layer_1_weights[27][30] + inp[31] * layer_1_weights[27][31] + inp[32] * layer_1_weights[27][32] + inp[33] * layer_1_weights[27][33] + inp[34] * layer_1_weights[27][34] + inp[35] * layer_1_weights[27][35] + inp[36] * layer_1_weights[27][36] + inp[37] * layer_1_weights[27][37] + inp[38] * layer_1_weights[27][38] + inp[39] * layer_1_weights[27][39] + inp[40] * layer_1_weights[27][40] + inp[41] * layer_1_weights[27][41] + inp[42] * layer_1_weights[27][42] + inp[43] * layer_1_weights[27][43] + inp[44] * layer_1_weights[27][44] + inp[45] * layer_1_weights[27][45] + inp[46] * layer_1_weights[27][46] + inp[47] * layer_1_weights[27][47] + inp[48] * layer_1_weights[27][48] + inp[49] * layer_1_weights[27][49] + inp[50] * layer_1_weights[27][50] + inp[51] * layer_1_weights[27][51] + inp[52] * layer_1_weights[27][52] + inp[53] * layer_1_weights[27][53] + inp[54] * layer_1_weights[27][54] + inp[55] * layer_1_weights[27][55] + inp[56] * layer_1_weights[27][56] + inp[57] * layer_1_weights[27][57] + inp[58] * layer_1_weights[27][58] + inp[59] * layer_1_weights[27][59] + inp[60] * layer_1_weights[27][60] + inp[61] * layer_1_weights[27][61] + inp[62] * layer_1_weights[27][62] + inp[63] * layer_1_weights[27][63] + inp[64] * layer_1_weights[27][64] + inp[65] * layer_1_weights[27][65] + inp[66] * layer_1_weights[27][66] + inp[67] * layer_1_weights[27][67] + inp[68] * layer_1_weights[27][68] + inp[69] * layer_1_weights[27][69] + inp[70] * layer_1_weights[27][70] + inp[71] * layer_1_weights[27][71] + inp[72] * layer_1_weights[27][72] + inp[73] * layer_1_weights[27][73] + inp[74] * layer_1_weights[27][74] + inp[75] * layer_1_weights[27][75] + inp[76] * layer_1_weights[27][76] + inp[77] * layer_1_weights[27][77] + inp[78] * layer_1_weights[27][78] + inp[79] * layer_1_weights[27][79] + inp[80] * layer_1_weights[27][80] + inp[81] * layer_1_weights[27][81] + inp[82] * layer_1_weights[27][82] + inp[83] * layer_1_weights[27][83] + inp[84] * layer_1_weights[27][84] + inp[85] * layer_1_weights[27][85] + inp[86] * layer_1_weights[27][86] + inp[87] * layer_1_weights[27][87] + inp[88] * layer_1_weights[27][88] + inp[89] * layer_1_weights[27][89] + inp[90] * layer_1_weights[27][90] + inp[91] * layer_1_weights[27][91] + inp[92] * layer_1_weights[27][92] + inp[93] * layer_1_weights[27][93] + inp[94] * layer_1_weights[27][94] + inp[95] * layer_1_weights[27][95] + inp[96] * layer_1_weights[27][96] + inp[97] * layer_1_weights[27][97] + inp[98] * layer_1_weights[27][98] + inp[99] * layer_1_weights[27][99] + inp[100] * layer_1_weights[27][100] + inp[101] * layer_1_weights[27][101] + inp[102] * layer_1_weights[27][102] + inp[103] * layer_1_weights[27][103] + inp[104] * layer_1_weights[27][104] + inp[105] * layer_1_weights[27][105] + inp[106] * layer_1_weights[27][106] + inp[107] * layer_1_weights[27][107] + inp[108] * layer_1_weights[27][108] + inp[109] * layer_1_weights[27][109] + inp[110] * layer_1_weights[27][110] + inp[111] * layer_1_weights[27][111] + inp[112] * layer_1_weights[27][112] + inp[113] * layer_1_weights[27][113] + inp[114] * layer_1_weights[27][114] + inp[115] * layer_1_weights[27][115] + inp[116] * layer_1_weights[27][116] + inp[117] * layer_1_weights[27][117] + inp[118] * layer_1_weights[27][118] + inp[119] * layer_1_weights[27][119] + inp[120] * layer_1_weights[27][120] + inp[121] * layer_1_weights[27][121] + inp[122] * layer_1_weights[27][122] + inp[123] * layer_1_weights[27][123] + inp[124] * layer_1_weights[27][124] + inp[125] * layer_1_weights[27][125] + inp[126] * layer_1_weights[27][126] + inp[127] * layer_1_weights[27][127] + inp[128] * layer_1_weights[27][128] + inp[129] * layer_1_weights[27][129] + inp[130] * layer_1_weights[27][130] + inp[131] * layer_1_weights[27][131] + inp[132] * layer_1_weights[27][132] + inp[133] * layer_1_weights[27][133] + inp[134] * layer_1_weights[27][134] + inp[135] * layer_1_weights[27][135] + inp[136] * layer_1_weights[27][136] + inp[137] * layer_1_weights[27][137] + inp[138] * layer_1_weights[27][138] + inp[139] * layer_1_weights[27][139] + inp[140] * layer_1_weights[27][140] + inp[141] * layer_1_weights[27][141] + inp[142] * layer_1_weights[27][142] + inp[143] * layer_1_weights[27][143]);
    assign layer_1_output_28 = relu(layer_1_biases[28] + inp[0] * layer_1_weights[28][0] + inp[1] * layer_1_weights[28][1] + inp[2] * layer_1_weights[28][2] + inp[3] * layer_1_weights[28][3] + inp[4] * layer_1_weights[28][4] + inp[5] * layer_1_weights[28][5] + inp[6] * layer_1_weights[28][6] + inp[7] * layer_1_weights[28][7] + inp[8] * layer_1_weights[28][8] + inp[9] * layer_1_weights[28][9] + inp[10] * layer_1_weights[28][10] + inp[11] * layer_1_weights[28][11] + inp[12] * layer_1_weights[28][12] + inp[13] * layer_1_weights[28][13] + inp[14] * layer_1_weights[28][14] + inp[15] * layer_1_weights[28][15] + inp[16] * layer_1_weights[28][16] + inp[17] * layer_1_weights[28][17] + inp[18] * layer_1_weights[28][18] + inp[19] * layer_1_weights[28][19] + inp[20] * layer_1_weights[28][20] + inp[21] * layer_1_weights[28][21] + inp[22] * layer_1_weights[28][22] + inp[23] * layer_1_weights[28][23] + inp[24] * layer_1_weights[28][24] + inp[25] * layer_1_weights[28][25] + inp[26] * layer_1_weights[28][26] + inp[27] * layer_1_weights[28][27] + inp[28] * layer_1_weights[28][28] + inp[29] * layer_1_weights[28][29] + inp[30] * layer_1_weights[28][30] + inp[31] * layer_1_weights[28][31] + inp[32] * layer_1_weights[28][32] + inp[33] * layer_1_weights[28][33] + inp[34] * layer_1_weights[28][34] + inp[35] * layer_1_weights[28][35] + inp[36] * layer_1_weights[28][36] + inp[37] * layer_1_weights[28][37] + inp[38] * layer_1_weights[28][38] + inp[39] * layer_1_weights[28][39] + inp[40] * layer_1_weights[28][40] + inp[41] * layer_1_weights[28][41] + inp[42] * layer_1_weights[28][42] + inp[43] * layer_1_weights[28][43] + inp[44] * layer_1_weights[28][44] + inp[45] * layer_1_weights[28][45] + inp[46] * layer_1_weights[28][46] + inp[47] * layer_1_weights[28][47] + inp[48] * layer_1_weights[28][48] + inp[49] * layer_1_weights[28][49] + inp[50] * layer_1_weights[28][50] + inp[51] * layer_1_weights[28][51] + inp[52] * layer_1_weights[28][52] + inp[53] * layer_1_weights[28][53] + inp[54] * layer_1_weights[28][54] + inp[55] * layer_1_weights[28][55] + inp[56] * layer_1_weights[28][56] + inp[57] * layer_1_weights[28][57] + inp[58] * layer_1_weights[28][58] + inp[59] * layer_1_weights[28][59] + inp[60] * layer_1_weights[28][60] + inp[61] * layer_1_weights[28][61] + inp[62] * layer_1_weights[28][62] + inp[63] * layer_1_weights[28][63] + inp[64] * layer_1_weights[28][64] + inp[65] * layer_1_weights[28][65] + inp[66] * layer_1_weights[28][66] + inp[67] * layer_1_weights[28][67] + inp[68] * layer_1_weights[28][68] + inp[69] * layer_1_weights[28][69] + inp[70] * layer_1_weights[28][70] + inp[71] * layer_1_weights[28][71] + inp[72] * layer_1_weights[28][72] + inp[73] * layer_1_weights[28][73] + inp[74] * layer_1_weights[28][74] + inp[75] * layer_1_weights[28][75] + inp[76] * layer_1_weights[28][76] + inp[77] * layer_1_weights[28][77] + inp[78] * layer_1_weights[28][78] + inp[79] * layer_1_weights[28][79] + inp[80] * layer_1_weights[28][80] + inp[81] * layer_1_weights[28][81] + inp[82] * layer_1_weights[28][82] + inp[83] * layer_1_weights[28][83] + inp[84] * layer_1_weights[28][84] + inp[85] * layer_1_weights[28][85] + inp[86] * layer_1_weights[28][86] + inp[87] * layer_1_weights[28][87] + inp[88] * layer_1_weights[28][88] + inp[89] * layer_1_weights[28][89] + inp[90] * layer_1_weights[28][90] + inp[91] * layer_1_weights[28][91] + inp[92] * layer_1_weights[28][92] + inp[93] * layer_1_weights[28][93] + inp[94] * layer_1_weights[28][94] + inp[95] * layer_1_weights[28][95] + inp[96] * layer_1_weights[28][96] + inp[97] * layer_1_weights[28][97] + inp[98] * layer_1_weights[28][98] + inp[99] * layer_1_weights[28][99] + inp[100] * layer_1_weights[28][100] + inp[101] * layer_1_weights[28][101] + inp[102] * layer_1_weights[28][102] + inp[103] * layer_1_weights[28][103] + inp[104] * layer_1_weights[28][104] + inp[105] * layer_1_weights[28][105] + inp[106] * layer_1_weights[28][106] + inp[107] * layer_1_weights[28][107] + inp[108] * layer_1_weights[28][108] + inp[109] * layer_1_weights[28][109] + inp[110] * layer_1_weights[28][110] + inp[111] * layer_1_weights[28][111] + inp[112] * layer_1_weights[28][112] + inp[113] * layer_1_weights[28][113] + inp[114] * layer_1_weights[28][114] + inp[115] * layer_1_weights[28][115] + inp[116] * layer_1_weights[28][116] + inp[117] * layer_1_weights[28][117] + inp[118] * layer_1_weights[28][118] + inp[119] * layer_1_weights[28][119] + inp[120] * layer_1_weights[28][120] + inp[121] * layer_1_weights[28][121] + inp[122] * layer_1_weights[28][122] + inp[123] * layer_1_weights[28][123] + inp[124] * layer_1_weights[28][124] + inp[125] * layer_1_weights[28][125] + inp[126] * layer_1_weights[28][126] + inp[127] * layer_1_weights[28][127] + inp[128] * layer_1_weights[28][128] + inp[129] * layer_1_weights[28][129] + inp[130] * layer_1_weights[28][130] + inp[131] * layer_1_weights[28][131] + inp[132] * layer_1_weights[28][132] + inp[133] * layer_1_weights[28][133] + inp[134] * layer_1_weights[28][134] + inp[135] * layer_1_weights[28][135] + inp[136] * layer_1_weights[28][136] + inp[137] * layer_1_weights[28][137] + inp[138] * layer_1_weights[28][138] + inp[139] * layer_1_weights[28][139] + inp[140] * layer_1_weights[28][140] + inp[141] * layer_1_weights[28][141] + inp[142] * layer_1_weights[28][142] + inp[143] * layer_1_weights[28][143]);
    assign layer_1_output_29 = relu(layer_1_biases[29] + inp[0] * layer_1_weights[29][0] + inp[1] * layer_1_weights[29][1] + inp[2] * layer_1_weights[29][2] + inp[3] * layer_1_weights[29][3] + inp[4] * layer_1_weights[29][4] + inp[5] * layer_1_weights[29][5] + inp[6] * layer_1_weights[29][6] + inp[7] * layer_1_weights[29][7] + inp[8] * layer_1_weights[29][8] + inp[9] * layer_1_weights[29][9] + inp[10] * layer_1_weights[29][10] + inp[11] * layer_1_weights[29][11] + inp[12] * layer_1_weights[29][12] + inp[13] * layer_1_weights[29][13] + inp[14] * layer_1_weights[29][14] + inp[15] * layer_1_weights[29][15] + inp[16] * layer_1_weights[29][16] + inp[17] * layer_1_weights[29][17] + inp[18] * layer_1_weights[29][18] + inp[19] * layer_1_weights[29][19] + inp[20] * layer_1_weights[29][20] + inp[21] * layer_1_weights[29][21] + inp[22] * layer_1_weights[29][22] + inp[23] * layer_1_weights[29][23] + inp[24] * layer_1_weights[29][24] + inp[25] * layer_1_weights[29][25] + inp[26] * layer_1_weights[29][26] + inp[27] * layer_1_weights[29][27] + inp[28] * layer_1_weights[29][28] + inp[29] * layer_1_weights[29][29] + inp[30] * layer_1_weights[29][30] + inp[31] * layer_1_weights[29][31] + inp[32] * layer_1_weights[29][32] + inp[33] * layer_1_weights[29][33] + inp[34] * layer_1_weights[29][34] + inp[35] * layer_1_weights[29][35] + inp[36] * layer_1_weights[29][36] + inp[37] * layer_1_weights[29][37] + inp[38] * layer_1_weights[29][38] + inp[39] * layer_1_weights[29][39] + inp[40] * layer_1_weights[29][40] + inp[41] * layer_1_weights[29][41] + inp[42] * layer_1_weights[29][42] + inp[43] * layer_1_weights[29][43] + inp[44] * layer_1_weights[29][44] + inp[45] * layer_1_weights[29][45] + inp[46] * layer_1_weights[29][46] + inp[47] * layer_1_weights[29][47] + inp[48] * layer_1_weights[29][48] + inp[49] * layer_1_weights[29][49] + inp[50] * layer_1_weights[29][50] + inp[51] * layer_1_weights[29][51] + inp[52] * layer_1_weights[29][52] + inp[53] * layer_1_weights[29][53] + inp[54] * layer_1_weights[29][54] + inp[55] * layer_1_weights[29][55] + inp[56] * layer_1_weights[29][56] + inp[57] * layer_1_weights[29][57] + inp[58] * layer_1_weights[29][58] + inp[59] * layer_1_weights[29][59] + inp[60] * layer_1_weights[29][60] + inp[61] * layer_1_weights[29][61] + inp[62] * layer_1_weights[29][62] + inp[63] * layer_1_weights[29][63] + inp[64] * layer_1_weights[29][64] + inp[65] * layer_1_weights[29][65] + inp[66] * layer_1_weights[29][66] + inp[67] * layer_1_weights[29][67] + inp[68] * layer_1_weights[29][68] + inp[69] * layer_1_weights[29][69] + inp[70] * layer_1_weights[29][70] + inp[71] * layer_1_weights[29][71] + inp[72] * layer_1_weights[29][72] + inp[73] * layer_1_weights[29][73] + inp[74] * layer_1_weights[29][74] + inp[75] * layer_1_weights[29][75] + inp[76] * layer_1_weights[29][76] + inp[77] * layer_1_weights[29][77] + inp[78] * layer_1_weights[29][78] + inp[79] * layer_1_weights[29][79] + inp[80] * layer_1_weights[29][80] + inp[81] * layer_1_weights[29][81] + inp[82] * layer_1_weights[29][82] + inp[83] * layer_1_weights[29][83] + inp[84] * layer_1_weights[29][84] + inp[85] * layer_1_weights[29][85] + inp[86] * layer_1_weights[29][86] + inp[87] * layer_1_weights[29][87] + inp[88] * layer_1_weights[29][88] + inp[89] * layer_1_weights[29][89] + inp[90] * layer_1_weights[29][90] + inp[91] * layer_1_weights[29][91] + inp[92] * layer_1_weights[29][92] + inp[93] * layer_1_weights[29][93] + inp[94] * layer_1_weights[29][94] + inp[95] * layer_1_weights[29][95] + inp[96] * layer_1_weights[29][96] + inp[97] * layer_1_weights[29][97] + inp[98] * layer_1_weights[29][98] + inp[99] * layer_1_weights[29][99] + inp[100] * layer_1_weights[29][100] + inp[101] * layer_1_weights[29][101] + inp[102] * layer_1_weights[29][102] + inp[103] * layer_1_weights[29][103] + inp[104] * layer_1_weights[29][104] + inp[105] * layer_1_weights[29][105] + inp[106] * layer_1_weights[29][106] + inp[107] * layer_1_weights[29][107] + inp[108] * layer_1_weights[29][108] + inp[109] * layer_1_weights[29][109] + inp[110] * layer_1_weights[29][110] + inp[111] * layer_1_weights[29][111] + inp[112] * layer_1_weights[29][112] + inp[113] * layer_1_weights[29][113] + inp[114] * layer_1_weights[29][114] + inp[115] * layer_1_weights[29][115] + inp[116] * layer_1_weights[29][116] + inp[117] * layer_1_weights[29][117] + inp[118] * layer_1_weights[29][118] + inp[119] * layer_1_weights[29][119] + inp[120] * layer_1_weights[29][120] + inp[121] * layer_1_weights[29][121] + inp[122] * layer_1_weights[29][122] + inp[123] * layer_1_weights[29][123] + inp[124] * layer_1_weights[29][124] + inp[125] * layer_1_weights[29][125] + inp[126] * layer_1_weights[29][126] + inp[127] * layer_1_weights[29][127] + inp[128] * layer_1_weights[29][128] + inp[129] * layer_1_weights[29][129] + inp[130] * layer_1_weights[29][130] + inp[131] * layer_1_weights[29][131] + inp[132] * layer_1_weights[29][132] + inp[133] * layer_1_weights[29][133] + inp[134] * layer_1_weights[29][134] + inp[135] * layer_1_weights[29][135] + inp[136] * layer_1_weights[29][136] + inp[137] * layer_1_weights[29][137] + inp[138] * layer_1_weights[29][138] + inp[139] * layer_1_weights[29][139] + inp[140] * layer_1_weights[29][140] + inp[141] * layer_1_weights[29][141] + inp[142] * layer_1_weights[29][142] + inp[143] * layer_1_weights[29][143]);
    assign layer_1_output_30 = relu(layer_1_biases[30] + inp[0] * layer_1_weights[30][0] + inp[1] * layer_1_weights[30][1] + inp[2] * layer_1_weights[30][2] + inp[3] * layer_1_weights[30][3] + inp[4] * layer_1_weights[30][4] + inp[5] * layer_1_weights[30][5] + inp[6] * layer_1_weights[30][6] + inp[7] * layer_1_weights[30][7] + inp[8] * layer_1_weights[30][8] + inp[9] * layer_1_weights[30][9] + inp[10] * layer_1_weights[30][10] + inp[11] * layer_1_weights[30][11] + inp[12] * layer_1_weights[30][12] + inp[13] * layer_1_weights[30][13] + inp[14] * layer_1_weights[30][14] + inp[15] * layer_1_weights[30][15] + inp[16] * layer_1_weights[30][16] + inp[17] * layer_1_weights[30][17] + inp[18] * layer_1_weights[30][18] + inp[19] * layer_1_weights[30][19] + inp[20] * layer_1_weights[30][20] + inp[21] * layer_1_weights[30][21] + inp[22] * layer_1_weights[30][22] + inp[23] * layer_1_weights[30][23] + inp[24] * layer_1_weights[30][24] + inp[25] * layer_1_weights[30][25] + inp[26] * layer_1_weights[30][26] + inp[27] * layer_1_weights[30][27] + inp[28] * layer_1_weights[30][28] + inp[29] * layer_1_weights[30][29] + inp[30] * layer_1_weights[30][30] + inp[31] * layer_1_weights[30][31] + inp[32] * layer_1_weights[30][32] + inp[33] * layer_1_weights[30][33] + inp[34] * layer_1_weights[30][34] + inp[35] * layer_1_weights[30][35] + inp[36] * layer_1_weights[30][36] + inp[37] * layer_1_weights[30][37] + inp[38] * layer_1_weights[30][38] + inp[39] * layer_1_weights[30][39] + inp[40] * layer_1_weights[30][40] + inp[41] * layer_1_weights[30][41] + inp[42] * layer_1_weights[30][42] + inp[43] * layer_1_weights[30][43] + inp[44] * layer_1_weights[30][44] + inp[45] * layer_1_weights[30][45] + inp[46] * layer_1_weights[30][46] + inp[47] * layer_1_weights[30][47] + inp[48] * layer_1_weights[30][48] + inp[49] * layer_1_weights[30][49] + inp[50] * layer_1_weights[30][50] + inp[51] * layer_1_weights[30][51] + inp[52] * layer_1_weights[30][52] + inp[53] * layer_1_weights[30][53] + inp[54] * layer_1_weights[30][54] + inp[55] * layer_1_weights[30][55] + inp[56] * layer_1_weights[30][56] + inp[57] * layer_1_weights[30][57] + inp[58] * layer_1_weights[30][58] + inp[59] * layer_1_weights[30][59] + inp[60] * layer_1_weights[30][60] + inp[61] * layer_1_weights[30][61] + inp[62] * layer_1_weights[30][62] + inp[63] * layer_1_weights[30][63] + inp[64] * layer_1_weights[30][64] + inp[65] * layer_1_weights[30][65] + inp[66] * layer_1_weights[30][66] + inp[67] * layer_1_weights[30][67] + inp[68] * layer_1_weights[30][68] + inp[69] * layer_1_weights[30][69] + inp[70] * layer_1_weights[30][70] + inp[71] * layer_1_weights[30][71] + inp[72] * layer_1_weights[30][72] + inp[73] * layer_1_weights[30][73] + inp[74] * layer_1_weights[30][74] + inp[75] * layer_1_weights[30][75] + inp[76] * layer_1_weights[30][76] + inp[77] * layer_1_weights[30][77] + inp[78] * layer_1_weights[30][78] + inp[79] * layer_1_weights[30][79] + inp[80] * layer_1_weights[30][80] + inp[81] * layer_1_weights[30][81] + inp[82] * layer_1_weights[30][82] + inp[83] * layer_1_weights[30][83] + inp[84] * layer_1_weights[30][84] + inp[85] * layer_1_weights[30][85] + inp[86] * layer_1_weights[30][86] + inp[87] * layer_1_weights[30][87] + inp[88] * layer_1_weights[30][88] + inp[89] * layer_1_weights[30][89] + inp[90] * layer_1_weights[30][90] + inp[91] * layer_1_weights[30][91] + inp[92] * layer_1_weights[30][92] + inp[93] * layer_1_weights[30][93] + inp[94] * layer_1_weights[30][94] + inp[95] * layer_1_weights[30][95] + inp[96] * layer_1_weights[30][96] + inp[97] * layer_1_weights[30][97] + inp[98] * layer_1_weights[30][98] + inp[99] * layer_1_weights[30][99] + inp[100] * layer_1_weights[30][100] + inp[101] * layer_1_weights[30][101] + inp[102] * layer_1_weights[30][102] + inp[103] * layer_1_weights[30][103] + inp[104] * layer_1_weights[30][104] + inp[105] * layer_1_weights[30][105] + inp[106] * layer_1_weights[30][106] + inp[107] * layer_1_weights[30][107] + inp[108] * layer_1_weights[30][108] + inp[109] * layer_1_weights[30][109] + inp[110] * layer_1_weights[30][110] + inp[111] * layer_1_weights[30][111] + inp[112] * layer_1_weights[30][112] + inp[113] * layer_1_weights[30][113] + inp[114] * layer_1_weights[30][114] + inp[115] * layer_1_weights[30][115] + inp[116] * layer_1_weights[30][116] + inp[117] * layer_1_weights[30][117] + inp[118] * layer_1_weights[30][118] + inp[119] * layer_1_weights[30][119] + inp[120] * layer_1_weights[30][120] + inp[121] * layer_1_weights[30][121] + inp[122] * layer_1_weights[30][122] + inp[123] * layer_1_weights[30][123] + inp[124] * layer_1_weights[30][124] + inp[125] * layer_1_weights[30][125] + inp[126] * layer_1_weights[30][126] + inp[127] * layer_1_weights[30][127] + inp[128] * layer_1_weights[30][128] + inp[129] * layer_1_weights[30][129] + inp[130] * layer_1_weights[30][130] + inp[131] * layer_1_weights[30][131] + inp[132] * layer_1_weights[30][132] + inp[133] * layer_1_weights[30][133] + inp[134] * layer_1_weights[30][134] + inp[135] * layer_1_weights[30][135] + inp[136] * layer_1_weights[30][136] + inp[137] * layer_1_weights[30][137] + inp[138] * layer_1_weights[30][138] + inp[139] * layer_1_weights[30][139] + inp[140] * layer_1_weights[30][140] + inp[141] * layer_1_weights[30][141] + inp[142] * layer_1_weights[30][142] + inp[143] * layer_1_weights[30][143]);
    assign layer_1_output_31 = relu(layer_1_biases[31] + inp[0] * layer_1_weights[31][0] + inp[1] * layer_1_weights[31][1] + inp[2] * layer_1_weights[31][2] + inp[3] * layer_1_weights[31][3] + inp[4] * layer_1_weights[31][4] + inp[5] * layer_1_weights[31][5] + inp[6] * layer_1_weights[31][6] + inp[7] * layer_1_weights[31][7] + inp[8] * layer_1_weights[31][8] + inp[9] * layer_1_weights[31][9] + inp[10] * layer_1_weights[31][10] + inp[11] * layer_1_weights[31][11] + inp[12] * layer_1_weights[31][12] + inp[13] * layer_1_weights[31][13] + inp[14] * layer_1_weights[31][14] + inp[15] * layer_1_weights[31][15] + inp[16] * layer_1_weights[31][16] + inp[17] * layer_1_weights[31][17] + inp[18] * layer_1_weights[31][18] + inp[19] * layer_1_weights[31][19] + inp[20] * layer_1_weights[31][20] + inp[21] * layer_1_weights[31][21] + inp[22] * layer_1_weights[31][22] + inp[23] * layer_1_weights[31][23] + inp[24] * layer_1_weights[31][24] + inp[25] * layer_1_weights[31][25] + inp[26] * layer_1_weights[31][26] + inp[27] * layer_1_weights[31][27] + inp[28] * layer_1_weights[31][28] + inp[29] * layer_1_weights[31][29] + inp[30] * layer_1_weights[31][30] + inp[31] * layer_1_weights[31][31] + inp[32] * layer_1_weights[31][32] + inp[33] * layer_1_weights[31][33] + inp[34] * layer_1_weights[31][34] + inp[35] * layer_1_weights[31][35] + inp[36] * layer_1_weights[31][36] + inp[37] * layer_1_weights[31][37] + inp[38] * layer_1_weights[31][38] + inp[39] * layer_1_weights[31][39] + inp[40] * layer_1_weights[31][40] + inp[41] * layer_1_weights[31][41] + inp[42] * layer_1_weights[31][42] + inp[43] * layer_1_weights[31][43] + inp[44] * layer_1_weights[31][44] + inp[45] * layer_1_weights[31][45] + inp[46] * layer_1_weights[31][46] + inp[47] * layer_1_weights[31][47] + inp[48] * layer_1_weights[31][48] + inp[49] * layer_1_weights[31][49] + inp[50] * layer_1_weights[31][50] + inp[51] * layer_1_weights[31][51] + inp[52] * layer_1_weights[31][52] + inp[53] * layer_1_weights[31][53] + inp[54] * layer_1_weights[31][54] + inp[55] * layer_1_weights[31][55] + inp[56] * layer_1_weights[31][56] + inp[57] * layer_1_weights[31][57] + inp[58] * layer_1_weights[31][58] + inp[59] * layer_1_weights[31][59] + inp[60] * layer_1_weights[31][60] + inp[61] * layer_1_weights[31][61] + inp[62] * layer_1_weights[31][62] + inp[63] * layer_1_weights[31][63] + inp[64] * layer_1_weights[31][64] + inp[65] * layer_1_weights[31][65] + inp[66] * layer_1_weights[31][66] + inp[67] * layer_1_weights[31][67] + inp[68] * layer_1_weights[31][68] + inp[69] * layer_1_weights[31][69] + inp[70] * layer_1_weights[31][70] + inp[71] * layer_1_weights[31][71] + inp[72] * layer_1_weights[31][72] + inp[73] * layer_1_weights[31][73] + inp[74] * layer_1_weights[31][74] + inp[75] * layer_1_weights[31][75] + inp[76] * layer_1_weights[31][76] + inp[77] * layer_1_weights[31][77] + inp[78] * layer_1_weights[31][78] + inp[79] * layer_1_weights[31][79] + inp[80] * layer_1_weights[31][80] + inp[81] * layer_1_weights[31][81] + inp[82] * layer_1_weights[31][82] + inp[83] * layer_1_weights[31][83] + inp[84] * layer_1_weights[31][84] + inp[85] * layer_1_weights[31][85] + inp[86] * layer_1_weights[31][86] + inp[87] * layer_1_weights[31][87] + inp[88] * layer_1_weights[31][88] + inp[89] * layer_1_weights[31][89] + inp[90] * layer_1_weights[31][90] + inp[91] * layer_1_weights[31][91] + inp[92] * layer_1_weights[31][92] + inp[93] * layer_1_weights[31][93] + inp[94] * layer_1_weights[31][94] + inp[95] * layer_1_weights[31][95] + inp[96] * layer_1_weights[31][96] + inp[97] * layer_1_weights[31][97] + inp[98] * layer_1_weights[31][98] + inp[99] * layer_1_weights[31][99] + inp[100] * layer_1_weights[31][100] + inp[101] * layer_1_weights[31][101] + inp[102] * layer_1_weights[31][102] + inp[103] * layer_1_weights[31][103] + inp[104] * layer_1_weights[31][104] + inp[105] * layer_1_weights[31][105] + inp[106] * layer_1_weights[31][106] + inp[107] * layer_1_weights[31][107] + inp[108] * layer_1_weights[31][108] + inp[109] * layer_1_weights[31][109] + inp[110] * layer_1_weights[31][110] + inp[111] * layer_1_weights[31][111] + inp[112] * layer_1_weights[31][112] + inp[113] * layer_1_weights[31][113] + inp[114] * layer_1_weights[31][114] + inp[115] * layer_1_weights[31][115] + inp[116] * layer_1_weights[31][116] + inp[117] * layer_1_weights[31][117] + inp[118] * layer_1_weights[31][118] + inp[119] * layer_1_weights[31][119] + inp[120] * layer_1_weights[31][120] + inp[121] * layer_1_weights[31][121] + inp[122] * layer_1_weights[31][122] + inp[123] * layer_1_weights[31][123] + inp[124] * layer_1_weights[31][124] + inp[125] * layer_1_weights[31][125] + inp[126] * layer_1_weights[31][126] + inp[127] * layer_1_weights[31][127] + inp[128] * layer_1_weights[31][128] + inp[129] * layer_1_weights[31][129] + inp[130] * layer_1_weights[31][130] + inp[131] * layer_1_weights[31][131] + inp[132] * layer_1_weights[31][132] + inp[133] * layer_1_weights[31][133] + inp[134] * layer_1_weights[31][134] + inp[135] * layer_1_weights[31][135] + inp[136] * layer_1_weights[31][136] + inp[137] * layer_1_weights[31][137] + inp[138] * layer_1_weights[31][138] + inp[139] * layer_1_weights[31][139] + inp[140] * layer_1_weights[31][140] + inp[141] * layer_1_weights[31][141] + inp[142] * layer_1_weights[31][142] + inp[143] * layer_1_weights[31][143]);

    // Layer 2: Dense
    wire signed [5:0] layer_2_weights [9:0][31:0];
    wire signed [5:0] layer_2_biases [9:0];

    assign layer_2_weights[0][0] = -6'sd7;
    assign layer_2_weights[0][1] = -6'sd11;
    assign layer_2_weights[0][2] = -6'sd3;
    assign layer_2_weights[0][3] = 6'sd1;
    assign layer_2_weights[0][4] = -6'sd16;
    assign layer_2_weights[0][5] = 6'sd4;
    assign layer_2_weights[0][6] = -6'sd12;
    assign layer_2_weights[0][7] = -6'sd4;
    assign layer_2_weights[0][8] = 6'sd7;
    assign layer_2_weights[0][9] = 6'sd2;
    assign layer_2_weights[0][10] = 6'sd5;
    assign layer_2_weights[0][11] = -6'sd3;
    assign layer_2_weights[0][12] = 6'sd7;
    assign layer_2_weights[0][13] = -6'sd10;
    assign layer_2_weights[0][14] = -6'sd2;
    assign layer_2_weights[0][15] = 6'sd5;
    assign layer_2_weights[0][16] = -6'sd6;
    assign layer_2_weights[0][17] = 6'sd9;
    assign layer_2_weights[0][18] = 6'sd14;
    assign layer_2_weights[0][19] = 6'sd1;
    assign layer_2_weights[0][20] = 6'sd2;
    assign layer_2_weights[0][21] = -6'sd8;
    assign layer_2_weights[0][22] = -6'sd11;
    assign layer_2_weights[0][23] = -6'sd13;
    assign layer_2_weights[0][24] = 6'sd6;
    assign layer_2_weights[0][25] = -6'sd6;
    assign layer_2_weights[0][26] = -6'sd4;
    assign layer_2_weights[0][27] = 6'sd0;
    assign layer_2_weights[0][28] = -6'sd5;
    assign layer_2_weights[0][29] = 6'sd0;
    assign layer_2_weights[0][30] = 6'sd6;
    assign layer_2_weights[0][31] = 6'sd4;
    assign layer_2_biases[0] = -6'sd6;
    assign layer_2_weights[1][0] = 6'sd6;
    assign layer_2_weights[1][1] = 6'sd8;
    assign layer_2_weights[1][2] = 6'sd3;
    assign layer_2_weights[1][3] = 6'sd7;
    assign layer_2_weights[1][4] = 6'sd4;
    assign layer_2_weights[1][5] = -6'sd11;
    assign layer_2_weights[1][6] = -6'sd7;
    assign layer_2_weights[1][7] = 6'sd1;
    assign layer_2_weights[1][8] = 6'sd3;
    assign layer_2_weights[1][9] = 6'sd9;
    assign layer_2_weights[1][10] = -6'sd10;
    assign layer_2_weights[1][11] = 6'sd7;
    assign layer_2_weights[1][12] = -6'sd6;
    assign layer_2_weights[1][13] = 6'sd0;
    assign layer_2_weights[1][14] = 6'sd1;
    assign layer_2_weights[1][15] = -6'sd9;
    assign layer_2_weights[1][16] = 6'sd5;
    assign layer_2_weights[1][17] = -6'sd14;
    assign layer_2_weights[1][18] = -6'sd9;
    assign layer_2_weights[1][19] = -6'sd9;
    assign layer_2_weights[1][20] = -6'sd10;
    assign layer_2_weights[1][21] = -6'sd3;
    assign layer_2_weights[1][22] = 6'sd1;
    assign layer_2_weights[1][23] = 6'sd5;
    assign layer_2_weights[1][24] = -6'sd4;
    assign layer_2_weights[1][25] = 6'sd5;
    assign layer_2_weights[1][26] = -6'sd4;
    assign layer_2_weights[1][27] = -6'sd18;
    assign layer_2_weights[1][28] = 6'sd5;
    assign layer_2_weights[1][29] = -6'sd11;
    assign layer_2_weights[1][30] = -6'sd10;
    assign layer_2_weights[1][31] = 6'sd5;
    assign layer_2_biases[1] = 6'sd5;
    assign layer_2_weights[2][0] = 6'sd8;
    assign layer_2_weights[2][1] = 6'sd0;
    assign layer_2_weights[2][2] = -6'sd16;
    assign layer_2_weights[2][3] = 6'sd8;
    assign layer_2_weights[2][4] = 6'sd6;
    assign layer_2_weights[2][5] = -6'sd1;
    assign layer_2_weights[2][6] = -6'sd5;
    assign layer_2_weights[2][7] = 6'sd8;
    assign layer_2_weights[2][8] = -6'sd3;
    assign layer_2_weights[2][9] = 6'sd6;
    assign layer_2_weights[2][10] = -6'sd16;
    assign layer_2_weights[2][11] = 6'sd6;
    assign layer_2_weights[2][12] = -6'sd11;
    assign layer_2_weights[2][13] = 6'sd6;
    assign layer_2_weights[2][14] = -6'sd2;
    assign layer_2_weights[2][15] = 6'sd9;
    assign layer_2_weights[2][16] = 6'sd6;
    assign layer_2_weights[2][17] = 6'sd13;
    assign layer_2_weights[2][18] = 6'sd3;
    assign layer_2_weights[2][19] = -6'sd1;
    assign layer_2_weights[2][20] = 6'sd3;
    assign layer_2_weights[2][21] = -6'sd5;
    assign layer_2_weights[2][22] = -6'sd3;
    assign layer_2_weights[2][23] = -6'sd10;
    assign layer_2_weights[2][24] = -6'sd2;
    assign layer_2_weights[2][25] = -6'sd16;
    assign layer_2_weights[2][26] = 6'sd0;
    assign layer_2_weights[2][27] = 6'sd0;
    assign layer_2_weights[2][28] = 6'sd7;
    assign layer_2_weights[2][29] = -6'sd1;
    assign layer_2_weights[2][30] = 6'sd1;
    assign layer_2_weights[2][31] = -6'sd9;
    assign layer_2_biases[2] = 6'sd1;
    assign layer_2_weights[3][0] = 6'sd5;
    assign layer_2_weights[3][1] = 6'sd8;
    assign layer_2_weights[3][2] = 6'sd3;
    assign layer_2_weights[3][3] = 6'sd4;
    assign layer_2_weights[3][4] = -6'sd13;
    assign layer_2_weights[3][5] = -6'sd7;
    assign layer_2_weights[3][6] = 6'sd2;
    assign layer_2_weights[3][7] = -6'sd2;
    assign layer_2_weights[3][8] = 6'sd3;
    assign layer_2_weights[3][9] = -6'sd6;
    assign layer_2_weights[3][10] = -6'sd4;
    assign layer_2_weights[3][11] = -6'sd2;
    assign layer_2_weights[3][12] = 6'sd5;
    assign layer_2_weights[3][13] = 6'sd6;
    assign layer_2_weights[3][14] = 6'sd0;
    assign layer_2_weights[3][15] = 6'sd1;
    assign layer_2_weights[3][16] = -6'sd4;
    assign layer_2_weights[3][17] = 6'sd5;
    assign layer_2_weights[3][18] = -6'sd9;
    assign layer_2_weights[3][19] = 6'sd4;
    assign layer_2_weights[3][20] = -6'sd7;
    assign layer_2_weights[3][21] = 6'sd4;
    assign layer_2_weights[3][22] = -6'sd1;
    assign layer_2_weights[3][23] = -6'sd14;
    assign layer_2_weights[3][24] = -6'sd13;
    assign layer_2_weights[3][25] = -6'sd9;
    assign layer_2_weights[3][26] = 6'sd6;
    assign layer_2_weights[3][27] = 6'sd0;
    assign layer_2_weights[3][28] = 6'sd0;
    assign layer_2_weights[3][29] = 6'sd4;
    assign layer_2_weights[3][30] = 6'sd4;
    assign layer_2_weights[3][31] = -6'sd1;
    assign layer_2_biases[3] = 6'sd0;
    assign layer_2_weights[4][0] = 6'sd7;
    assign layer_2_weights[4][1] = -6'sd6;
    assign layer_2_weights[4][2] = 6'sd7;
    assign layer_2_weights[4][3] = -6'sd5;
    assign layer_2_weights[4][4] = 6'sd6;
    assign layer_2_weights[4][5] = 6'sd1;
    assign layer_2_weights[4][6] = 6'sd5;
    assign layer_2_weights[4][7] = 6'sd5;
    assign layer_2_weights[4][8] = 6'sd0;
    assign layer_2_weights[4][9] = -6'sd6;
    assign layer_2_weights[4][10] = 6'sd1;
    assign layer_2_weights[4][11] = -6'sd6;
    assign layer_2_weights[4][12] = -6'sd6;
    assign layer_2_weights[4][13] = -6'sd5;
    assign layer_2_weights[4][14] = 6'sd13;
    assign layer_2_weights[4][15] = -6'sd16;
    assign layer_2_weights[4][16] = -6'sd6;
    assign layer_2_weights[4][17] = -6'sd14;
    assign layer_2_weights[4][18] = -6'sd1;
    assign layer_2_weights[4][19] = -6'sd14;
    assign layer_2_weights[4][20] = -6'sd4;
    assign layer_2_weights[4][21] = -6'sd15;
    assign layer_2_weights[4][22] = 6'sd6;
    assign layer_2_weights[4][23] = 6'sd5;
    assign layer_2_weights[4][24] = 6'sd7;
    assign layer_2_weights[4][25] = -6'sd14;
    assign layer_2_weights[4][26] = 6'sd2;
    assign layer_2_weights[4][27] = 6'sd6;
    assign layer_2_weights[4][28] = 6'sd2;
    assign layer_2_weights[4][29] = -6'sd10;
    assign layer_2_weights[4][30] = 6'sd0;
    assign layer_2_weights[4][31] = 6'sd5;
    assign layer_2_biases[4] = 6'sd3;
    assign layer_2_weights[5][0] = -6'sd2;
    assign layer_2_weights[5][1] = 6'sd6;
    assign layer_2_weights[5][2] = -6'sd4;
    assign layer_2_weights[5][3] = -6'sd14;
    assign layer_2_weights[5][4] = -6'sd6;
    assign layer_2_weights[5][5] = -6'sd6;
    assign layer_2_weights[5][6] = 6'sd9;
    assign layer_2_weights[5][7] = -6'sd5;
    assign layer_2_weights[5][8] = 6'sd3;
    assign layer_2_weights[5][9] = 6'sd2;
    assign layer_2_weights[5][10] = 6'sd3;
    assign layer_2_weights[5][11] = -6'sd5;
    assign layer_2_weights[5][12] = 6'sd7;
    assign layer_2_weights[5][13] = -6'sd4;
    assign layer_2_weights[5][14] = 6'sd3;
    assign layer_2_weights[5][15] = 6'sd1;
    assign layer_2_weights[5][16] = 6'sd3;
    assign layer_2_weights[5][17] = 6'sd1;
    assign layer_2_weights[5][18] = -6'sd17;
    assign layer_2_weights[5][19] = 6'sd7;
    assign layer_2_weights[5][20] = 6'sd0;
    assign layer_2_weights[5][21] = 6'sd12;
    assign layer_2_weights[5][22] = 6'sd0;
    assign layer_2_weights[5][23] = 6'sd2;
    assign layer_2_weights[5][24] = -6'sd2;
    assign layer_2_weights[5][25] = 6'sd17;
    assign layer_2_weights[5][26] = 6'sd0;
    assign layer_2_weights[5][27] = 6'sd2;
    assign layer_2_weights[5][28] = -6'sd9;
    assign layer_2_weights[5][29] = 6'sd5;
    assign layer_2_weights[5][30] = -6'sd6;
    assign layer_2_weights[5][31] = -6'sd10;
    assign layer_2_biases[5] = 6'sd2;
    assign layer_2_weights[6][0] = -6'sd10;
    assign layer_2_weights[6][1] = -6'sd15;
    assign layer_2_weights[6][2] = -6'sd2;
    assign layer_2_weights[6][3] = -6'sd13;
    assign layer_2_weights[6][4] = -6'sd2;
    assign layer_2_weights[6][5] = -6'sd1;
    assign layer_2_weights[6][6] = -6'sd11;
    assign layer_2_weights[6][7] = 6'sd5;
    assign layer_2_weights[6][8] = 6'sd4;
    assign layer_2_weights[6][9] = 6'sd3;
    assign layer_2_weights[6][10] = 6'sd6;
    assign layer_2_weights[6][11] = 6'sd0;
    assign layer_2_weights[6][12] = 6'sd7;
    assign layer_2_weights[6][13] = -6'sd16;
    assign layer_2_weights[6][14] = 6'sd2;
    assign layer_2_weights[6][15] = -6'sd8;
    assign layer_2_weights[6][16] = 6'sd6;
    assign layer_2_weights[6][17] = -6'sd8;
    assign layer_2_weights[6][18] = 6'sd2;
    assign layer_2_weights[6][19] = -6'sd6;
    assign layer_2_weights[6][20] = 6'sd2;
    assign layer_2_weights[6][21] = 6'sd7;
    assign layer_2_weights[6][22] = -6'sd1;
    assign layer_2_weights[6][23] = 6'sd2;
    assign layer_2_weights[6][24] = 6'sd3;
    assign layer_2_weights[6][25] = 6'sd2;
    assign layer_2_weights[6][26] = -6'sd15;
    assign layer_2_weights[6][27] = 6'sd4;
    assign layer_2_weights[6][28] = -6'sd1;
    assign layer_2_weights[6][29] = 6'sd8;
    assign layer_2_weights[6][30] = 6'sd1;
    assign layer_2_weights[6][31] = -6'sd9;
    assign layer_2_biases[6] = -6'sd1;
    assign layer_2_weights[7][0] = -6'sd8;
    assign layer_2_weights[7][1] = -6'sd8;
    assign layer_2_weights[7][2] = 6'sd0;
    assign layer_2_weights[7][3] = 6'sd2;
    assign layer_2_weights[7][4] = 6'sd7;
    assign layer_2_weights[7][5] = 6'sd4;
    assign layer_2_weights[7][6] = -6'sd4;
    assign layer_2_weights[7][7] = 6'sd1;
    assign layer_2_weights[7][8] = -6'sd5;
    assign layer_2_weights[7][9] = 6'sd5;
    assign layer_2_weights[7][10] = 6'sd2;
    assign layer_2_weights[7][11] = -6'sd11;
    assign layer_2_weights[7][12] = -6'sd10;
    assign layer_2_weights[7][13] = 6'sd7;
    assign layer_2_weights[7][14] = 6'sd0;
    assign layer_2_weights[7][15] = 6'sd6;
    assign layer_2_weights[7][16] = 6'sd6;
    assign layer_2_weights[7][17] = -6'sd5;
    assign layer_2_weights[7][18] = -6'sd1;
    assign layer_2_weights[7][19] = 6'sd6;
    assign layer_2_weights[7][20] = -6'sd8;
    assign layer_2_weights[7][21] = -6'sd10;
    assign layer_2_weights[7][22] = 6'sd4;
    assign layer_2_weights[7][23] = 6'sd0;
    assign layer_2_weights[7][24] = -6'sd10;
    assign layer_2_weights[7][25] = -6'sd2;
    assign layer_2_weights[7][26] = 6'sd6;
    assign layer_2_weights[7][27] = 6'sd4;
    assign layer_2_weights[7][28] = 6'sd3;
    assign layer_2_weights[7][29] = -6'sd13;
    assign layer_2_weights[7][30] = -6'sd4;
    assign layer_2_weights[7][31] = 6'sd9;
    assign layer_2_biases[7] = 6'sd4;
    assign layer_2_weights[8][0] = -6'sd8;
    assign layer_2_weights[8][1] = -6'sd6;
    assign layer_2_weights[8][2] = -6'sd14;
    assign layer_2_weights[8][3] = -6'sd2;
    assign layer_2_weights[8][4] = 6'sd9;
    assign layer_2_weights[8][5] = -6'sd15;
    assign layer_2_weights[8][6] = 6'sd4;
    assign layer_2_weights[8][7] = -6'sd15;
    assign layer_2_weights[8][8] = 6'sd7;
    assign layer_2_weights[8][9] = -6'sd11;
    assign layer_2_weights[8][10] = -6'sd8;
    assign layer_2_weights[8][11] = 6'sd2;
    assign layer_2_weights[8][12] = 6'sd5;
    assign layer_2_weights[8][13] = 6'sd6;
    assign layer_2_weights[8][14] = 6'sd1;
    assign layer_2_weights[8][15] = 6'sd0;
    assign layer_2_weights[8][16] = -6'sd1;
    assign layer_2_weights[8][17] = 6'sd8;
    assign layer_2_weights[8][18] = 6'sd0;
    assign layer_2_weights[8][19] = -6'sd4;
    assign layer_2_weights[8][20] = 6'sd3;
    assign layer_2_weights[8][21] = -6'sd1;
    assign layer_2_weights[8][22] = 6'sd4;
    assign layer_2_weights[8][23] = -6'sd1;
    assign layer_2_weights[8][24] = 6'sd1;
    assign layer_2_weights[8][25] = -6'sd3;
    assign layer_2_weights[8][26] = 6'sd2;
    assign layer_2_weights[8][27] = 6'sd5;
    assign layer_2_weights[8][28] = 6'sd5;
    assign layer_2_weights[8][29] = 6'sd1;
    assign layer_2_weights[8][30] = 6'sd0;
    assign layer_2_weights[8][31] = -6'sd1;
    assign layer_2_biases[8] = -6'sd4;
    assign layer_2_weights[9][0] = 6'sd2;
    assign layer_2_weights[9][1] = 6'sd12;
    assign layer_2_weights[9][2] = 6'sd9;
    assign layer_2_weights[9][3] = 6'sd4;
    assign layer_2_weights[9][4] = -6'sd4;
    assign layer_2_weights[9][5] = 6'sd8;
    assign layer_2_weights[9][6] = 6'sd4;
    assign layer_2_weights[9][7] = -6'sd10;
    assign layer_2_weights[9][8] = -6'sd3;
    assign layer_2_weights[9][9] = -6'sd11;
    assign layer_2_weights[9][10] = 6'sd2;
    assign layer_2_weights[9][11] = 6'sd2;
    assign layer_2_weights[9][12] = 6'sd1;
    assign layer_2_weights[9][13] = -6'sd15;
    assign layer_2_weights[9][14] = -6'sd14;
    assign layer_2_weights[9][15] = 6'sd1;
    assign layer_2_weights[9][16] = -6'sd21;
    assign layer_2_weights[9][17] = -6'sd10;
    assign layer_2_weights[9][18] = 6'sd3;
    assign layer_2_weights[9][19] = 6'sd3;
    assign layer_2_weights[9][20] = 6'sd5;
    assign layer_2_weights[9][21] = -6'sd2;
    assign layer_2_weights[9][22] = 6'sd4;
    assign layer_2_weights[9][23] = 6'sd4;
    assign layer_2_weights[9][24] = -6'sd5;
    assign layer_2_weights[9][25] = 6'sd1;
    assign layer_2_weights[9][26] = 6'sd4;
    assign layer_2_weights[9][27] = -6'sd6;
    assign layer_2_weights[9][28] = -6'sd12;
    assign layer_2_weights[9][29] = -6'sd21;
    assign layer_2_weights[9][30] = 6'sd4;
    assign layer_2_weights[9][31] = 6'sd4;
    assign layer_2_biases[9] = -6'sd2;

    wire signed [5:0] layer_2_output_0;
    wire signed [5:0] layer_2_output_1;
    wire signed [5:0] layer_2_output_2;
    wire signed [5:0] layer_2_output_3;
    wire signed [5:0] layer_2_output_4;
    wire signed [5:0] layer_2_output_5;
    wire signed [5:0] layer_2_output_6;
    wire signed [5:0] layer_2_output_7;
    wire signed [5:0] layer_2_output_8;
    wire signed [5:0] layer_2_output_9;
    assign layer_2_output_0 = relu(layer_2_biases[0] + inp[0] * layer_2_weights[0][0] + inp[1] * layer_2_weights[0][1] + inp[2] * layer_2_weights[0][2] + inp[3] * layer_2_weights[0][3] + inp[4] * layer_2_weights[0][4] + inp[5] * layer_2_weights[0][5] + inp[6] * layer_2_weights[0][6] + inp[7] * layer_2_weights[0][7] + inp[8] * layer_2_weights[0][8] + inp[9] * layer_2_weights[0][9] + inp[10] * layer_2_weights[0][10] + inp[11] * layer_2_weights[0][11] + inp[12] * layer_2_weights[0][12] + inp[13] * layer_2_weights[0][13] + inp[14] * layer_2_weights[0][14] + inp[15] * layer_2_weights[0][15] + inp[16] * layer_2_weights[0][16] + inp[17] * layer_2_weights[0][17] + inp[18] * layer_2_weights[0][18] + inp[19] * layer_2_weights[0][19] + inp[20] * layer_2_weights[0][20] + inp[21] * layer_2_weights[0][21] + inp[22] * layer_2_weights[0][22] + inp[23] * layer_2_weights[0][23] + inp[24] * layer_2_weights[0][24] + inp[25] * layer_2_weights[0][25] + inp[26] * layer_2_weights[0][26] + inp[27] * layer_2_weights[0][27] + inp[28] * layer_2_weights[0][28] + inp[29] * layer_2_weights[0][29] + inp[30] * layer_2_weights[0][30] + inp[31] * layer_2_weights[0][31]);
    assign layer_2_output_1 = relu(layer_2_biases[1] + inp[0] * layer_2_weights[1][0] + inp[1] * layer_2_weights[1][1] + inp[2] * layer_2_weights[1][2] + inp[3] * layer_2_weights[1][3] + inp[4] * layer_2_weights[1][4] + inp[5] * layer_2_weights[1][5] + inp[6] * layer_2_weights[1][6] + inp[7] * layer_2_weights[1][7] + inp[8] * layer_2_weights[1][8] + inp[9] * layer_2_weights[1][9] + inp[10] * layer_2_weights[1][10] + inp[11] * layer_2_weights[1][11] + inp[12] * layer_2_weights[1][12] + inp[13] * layer_2_weights[1][13] + inp[14] * layer_2_weights[1][14] + inp[15] * layer_2_weights[1][15] + inp[16] * layer_2_weights[1][16] + inp[17] * layer_2_weights[1][17] + inp[18] * layer_2_weights[1][18] + inp[19] * layer_2_weights[1][19] + inp[20] * layer_2_weights[1][20] + inp[21] * layer_2_weights[1][21] + inp[22] * layer_2_weights[1][22] + inp[23] * layer_2_weights[1][23] + inp[24] * layer_2_weights[1][24] + inp[25] * layer_2_weights[1][25] + inp[26] * layer_2_weights[1][26] + inp[27] * layer_2_weights[1][27] + inp[28] * layer_2_weights[1][28] + inp[29] * layer_2_weights[1][29] + inp[30] * layer_2_weights[1][30] + inp[31] * layer_2_weights[1][31]);
    assign layer_2_output_2 = relu(layer_2_biases[2] + inp[0] * layer_2_weights[2][0] + inp[1] * layer_2_weights[2][1] + inp[2] * layer_2_weights[2][2] + inp[3] * layer_2_weights[2][3] + inp[4] * layer_2_weights[2][4] + inp[5] * layer_2_weights[2][5] + inp[6] * layer_2_weights[2][6] + inp[7] * layer_2_weights[2][7] + inp[8] * layer_2_weights[2][8] + inp[9] * layer_2_weights[2][9] + inp[10] * layer_2_weights[2][10] + inp[11] * layer_2_weights[2][11] + inp[12] * layer_2_weights[2][12] + inp[13] * layer_2_weights[2][13] + inp[14] * layer_2_weights[2][14] + inp[15] * layer_2_weights[2][15] + inp[16] * layer_2_weights[2][16] + inp[17] * layer_2_weights[2][17] + inp[18] * layer_2_weights[2][18] + inp[19] * layer_2_weights[2][19] + inp[20] * layer_2_weights[2][20] + inp[21] * layer_2_weights[2][21] + inp[22] * layer_2_weights[2][22] + inp[23] * layer_2_weights[2][23] + inp[24] * layer_2_weights[2][24] + inp[25] * layer_2_weights[2][25] + inp[26] * layer_2_weights[2][26] + inp[27] * layer_2_weights[2][27] + inp[28] * layer_2_weights[2][28] + inp[29] * layer_2_weights[2][29] + inp[30] * layer_2_weights[2][30] + inp[31] * layer_2_weights[2][31]);
    assign layer_2_output_3 = relu(layer_2_biases[3] + inp[0] * layer_2_weights[3][0] + inp[1] * layer_2_weights[3][1] + inp[2] * layer_2_weights[3][2] + inp[3] * layer_2_weights[3][3] + inp[4] * layer_2_weights[3][4] + inp[5] * layer_2_weights[3][5] + inp[6] * layer_2_weights[3][6] + inp[7] * layer_2_weights[3][7] + inp[8] * layer_2_weights[3][8] + inp[9] * layer_2_weights[3][9] + inp[10] * layer_2_weights[3][10] + inp[11] * layer_2_weights[3][11] + inp[12] * layer_2_weights[3][12] + inp[13] * layer_2_weights[3][13] + inp[14] * layer_2_weights[3][14] + inp[15] * layer_2_weights[3][15] + inp[16] * layer_2_weights[3][16] + inp[17] * layer_2_weights[3][17] + inp[18] * layer_2_weights[3][18] + inp[19] * layer_2_weights[3][19] + inp[20] * layer_2_weights[3][20] + inp[21] * layer_2_weights[3][21] + inp[22] * layer_2_weights[3][22] + inp[23] * layer_2_weights[3][23] + inp[24] * layer_2_weights[3][24] + inp[25] * layer_2_weights[3][25] + inp[26] * layer_2_weights[3][26] + inp[27] * layer_2_weights[3][27] + inp[28] * layer_2_weights[3][28] + inp[29] * layer_2_weights[3][29] + inp[30] * layer_2_weights[3][30] + inp[31] * layer_2_weights[3][31]);
    assign layer_2_output_4 = relu(layer_2_biases[4] + inp[0] * layer_2_weights[4][0] + inp[1] * layer_2_weights[4][1] + inp[2] * layer_2_weights[4][2] + inp[3] * layer_2_weights[4][3] + inp[4] * layer_2_weights[4][4] + inp[5] * layer_2_weights[4][5] + inp[6] * layer_2_weights[4][6] + inp[7] * layer_2_weights[4][7] + inp[8] * layer_2_weights[4][8] + inp[9] * layer_2_weights[4][9] + inp[10] * layer_2_weights[4][10] + inp[11] * layer_2_weights[4][11] + inp[12] * layer_2_weights[4][12] + inp[13] * layer_2_weights[4][13] + inp[14] * layer_2_weights[4][14] + inp[15] * layer_2_weights[4][15] + inp[16] * layer_2_weights[4][16] + inp[17] * layer_2_weights[4][17] + inp[18] * layer_2_weights[4][18] + inp[19] * layer_2_weights[4][19] + inp[20] * layer_2_weights[4][20] + inp[21] * layer_2_weights[4][21] + inp[22] * layer_2_weights[4][22] + inp[23] * layer_2_weights[4][23] + inp[24] * layer_2_weights[4][24] + inp[25] * layer_2_weights[4][25] + inp[26] * layer_2_weights[4][26] + inp[27] * layer_2_weights[4][27] + inp[28] * layer_2_weights[4][28] + inp[29] * layer_2_weights[4][29] + inp[30] * layer_2_weights[4][30] + inp[31] * layer_2_weights[4][31]);
    assign layer_2_output_5 = relu(layer_2_biases[5] + inp[0] * layer_2_weights[5][0] + inp[1] * layer_2_weights[5][1] + inp[2] * layer_2_weights[5][2] + inp[3] * layer_2_weights[5][3] + inp[4] * layer_2_weights[5][4] + inp[5] * layer_2_weights[5][5] + inp[6] * layer_2_weights[5][6] + inp[7] * layer_2_weights[5][7] + inp[8] * layer_2_weights[5][8] + inp[9] * layer_2_weights[5][9] + inp[10] * layer_2_weights[5][10] + inp[11] * layer_2_weights[5][11] + inp[12] * layer_2_weights[5][12] + inp[13] * layer_2_weights[5][13] + inp[14] * layer_2_weights[5][14] + inp[15] * layer_2_weights[5][15] + inp[16] * layer_2_weights[5][16] + inp[17] * layer_2_weights[5][17] + inp[18] * layer_2_weights[5][18] + inp[19] * layer_2_weights[5][19] + inp[20] * layer_2_weights[5][20] + inp[21] * layer_2_weights[5][21] + inp[22] * layer_2_weights[5][22] + inp[23] * layer_2_weights[5][23] + inp[24] * layer_2_weights[5][24] + inp[25] * layer_2_weights[5][25] + inp[26] * layer_2_weights[5][26] + inp[27] * layer_2_weights[5][27] + inp[28] * layer_2_weights[5][28] + inp[29] * layer_2_weights[5][29] + inp[30] * layer_2_weights[5][30] + inp[31] * layer_2_weights[5][31]);
    assign layer_2_output_6 = relu(layer_2_biases[6] + inp[0] * layer_2_weights[6][0] + inp[1] * layer_2_weights[6][1] + inp[2] * layer_2_weights[6][2] + inp[3] * layer_2_weights[6][3] + inp[4] * layer_2_weights[6][4] + inp[5] * layer_2_weights[6][5] + inp[6] * layer_2_weights[6][6] + inp[7] * layer_2_weights[6][7] + inp[8] * layer_2_weights[6][8] + inp[9] * layer_2_weights[6][9] + inp[10] * layer_2_weights[6][10] + inp[11] * layer_2_weights[6][11] + inp[12] * layer_2_weights[6][12] + inp[13] * layer_2_weights[6][13] + inp[14] * layer_2_weights[6][14] + inp[15] * layer_2_weights[6][15] + inp[16] * layer_2_weights[6][16] + inp[17] * layer_2_weights[6][17] + inp[18] * layer_2_weights[6][18] + inp[19] * layer_2_weights[6][19] + inp[20] * layer_2_weights[6][20] + inp[21] * layer_2_weights[6][21] + inp[22] * layer_2_weights[6][22] + inp[23] * layer_2_weights[6][23] + inp[24] * layer_2_weights[6][24] + inp[25] * layer_2_weights[6][25] + inp[26] * layer_2_weights[6][26] + inp[27] * layer_2_weights[6][27] + inp[28] * layer_2_weights[6][28] + inp[29] * layer_2_weights[6][29] + inp[30] * layer_2_weights[6][30] + inp[31] * layer_2_weights[6][31]);
    assign layer_2_output_7 = relu(layer_2_biases[7] + inp[0] * layer_2_weights[7][0] + inp[1] * layer_2_weights[7][1] + inp[2] * layer_2_weights[7][2] + inp[3] * layer_2_weights[7][3] + inp[4] * layer_2_weights[7][4] + inp[5] * layer_2_weights[7][5] + inp[6] * layer_2_weights[7][6] + inp[7] * layer_2_weights[7][7] + inp[8] * layer_2_weights[7][8] + inp[9] * layer_2_weights[7][9] + inp[10] * layer_2_weights[7][10] + inp[11] * layer_2_weights[7][11] + inp[12] * layer_2_weights[7][12] + inp[13] * layer_2_weights[7][13] + inp[14] * layer_2_weights[7][14] + inp[15] * layer_2_weights[7][15] + inp[16] * layer_2_weights[7][16] + inp[17] * layer_2_weights[7][17] + inp[18] * layer_2_weights[7][18] + inp[19] * layer_2_weights[7][19] + inp[20] * layer_2_weights[7][20] + inp[21] * layer_2_weights[7][21] + inp[22] * layer_2_weights[7][22] + inp[23] * layer_2_weights[7][23] + inp[24] * layer_2_weights[7][24] + inp[25] * layer_2_weights[7][25] + inp[26] * layer_2_weights[7][26] + inp[27] * layer_2_weights[7][27] + inp[28] * layer_2_weights[7][28] + inp[29] * layer_2_weights[7][29] + inp[30] * layer_2_weights[7][30] + inp[31] * layer_2_weights[7][31]);
    assign layer_2_output_8 = relu(layer_2_biases[8] + inp[0] * layer_2_weights[8][0] + inp[1] * layer_2_weights[8][1] + inp[2] * layer_2_weights[8][2] + inp[3] * layer_2_weights[8][3] + inp[4] * layer_2_weights[8][4] + inp[5] * layer_2_weights[8][5] + inp[6] * layer_2_weights[8][6] + inp[7] * layer_2_weights[8][7] + inp[8] * layer_2_weights[8][8] + inp[9] * layer_2_weights[8][9] + inp[10] * layer_2_weights[8][10] + inp[11] * layer_2_weights[8][11] + inp[12] * layer_2_weights[8][12] + inp[13] * layer_2_weights[8][13] + inp[14] * layer_2_weights[8][14] + inp[15] * layer_2_weights[8][15] + inp[16] * layer_2_weights[8][16] + inp[17] * layer_2_weights[8][17] + inp[18] * layer_2_weights[8][18] + inp[19] * layer_2_weights[8][19] + inp[20] * layer_2_weights[8][20] + inp[21] * layer_2_weights[8][21] + inp[22] * layer_2_weights[8][22] + inp[23] * layer_2_weights[8][23] + inp[24] * layer_2_weights[8][24] + inp[25] * layer_2_weights[8][25] + inp[26] * layer_2_weights[8][26] + inp[27] * layer_2_weights[8][27] + inp[28] * layer_2_weights[8][28] + inp[29] * layer_2_weights[8][29] + inp[30] * layer_2_weights[8][30] + inp[31] * layer_2_weights[8][31]);
    assign layer_2_output_9 = relu(layer_2_biases[9] + inp[0] * layer_2_weights[9][0] + inp[1] * layer_2_weights[9][1] + inp[2] * layer_2_weights[9][2] + inp[3] * layer_2_weights[9][3] + inp[4] * layer_2_weights[9][4] + inp[5] * layer_2_weights[9][5] + inp[6] * layer_2_weights[9][6] + inp[7] * layer_2_weights[9][7] + inp[8] * layer_2_weights[9][8] + inp[9] * layer_2_weights[9][9] + inp[10] * layer_2_weights[9][10] + inp[11] * layer_2_weights[9][11] + inp[12] * layer_2_weights[9][12] + inp[13] * layer_2_weights[9][13] + inp[14] * layer_2_weights[9][14] + inp[15] * layer_2_weights[9][15] + inp[16] * layer_2_weights[9][16] + inp[17] * layer_2_weights[9][17] + inp[18] * layer_2_weights[9][18] + inp[19] * layer_2_weights[9][19] + inp[20] * layer_2_weights[9][20] + inp[21] * layer_2_weights[9][21] + inp[22] * layer_2_weights[9][22] + inp[23] * layer_2_weights[9][23] + inp[24] * layer_2_weights[9][24] + inp[25] * layer_2_weights[9][25] + inp[26] * layer_2_weights[9][26] + inp[27] * layer_2_weights[9][27] + inp[28] * layer_2_weights[9][28] + inp[29] * layer_2_weights[9][29] + inp[30] * layer_2_weights[9][30] + inp[31] * layer_2_weights[9][31]);

    // Softmax approximation: Winner-takes-all
    assign class = find_max(layer_2_output_0, layer_2_output_1, layer_2_output_2, layer_2_output_3, layer_2_output_4, layer_2_output_5, layer_2_output_6, layer_2_output_7, layer_2_output_8, layer_2_output_9);


    // ReLU function
    function signed [5:0] relu;
        input signed [5:0] x;
        begin
            if (x > 0)
                relu = x;
            else
                relu = 0;
        end
    endfunction

    // Find maximum value function
    function [3:0] find_max;
        input signed [5:0] out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9;
        integer i;
        reg signed [5:0] max_val;
        reg [3:0] max_idx;

        begin
            max_val = out_0;
            max_idx = 0;
            if (out_1 > max_val) begin
                max_val = out_1;
                max_idx = 1;
            end
            if (out_2 > max_val) begin
                max_val = out_2;
                max_idx = 2;
            end
            if (out_3 > max_val) begin
                max_val = out_3;
                max_idx = 3;
            end
            if (out_4 > max_val) begin
                max_val = out_4;
                max_idx = 4;
            end
            if (out_5 > max_val) begin
                max_val = out_5;
                max_idx = 5;
            end
            if (out_6 > max_val) begin
                max_val = out_6;
                max_idx = 6;
            end
            if (out_7 > max_val) begin
                max_val = out_7;
                max_idx = 7;
            end
            if (out_8 > max_val) begin
                max_val = out_8;
                max_idx = 8;
            end
            if (out_9 > max_val) begin
                max_val = out_9;
                max_idx = 9;
            end
            find_max = max_idx;
        end
    endfunction
endmodule
