module MLP_model (
    input predict,
    input [143:0] inp,
    output reg [3:0] class
);

    // Layer 1: Dense
    reg signed [7:0] layer_1_weights [143:0][7:0];
    reg signed [7:0] layer_1_biases [7:0];
    reg signed [15:0] layer_1_outputs [7:0];

    // Layer 2: Dense
    reg signed [7:0] layer_2_weights [7:0][9:0];
    reg signed [7:0] layer_2_biases [9:0];
    reg signed [23:0] layer_2_outputs [9:0];

    reg signed [23:0] max_val;
    reg [3:0] max_idx;

    initial begin
        layer_1_weights[0][0] = 3;
        layer_1_weights[1][0] = -2;
        layer_1_weights[2][0] = 19;
        layer_1_weights[3][0] = 20;
        layer_1_weights[4][0] = 8;
        layer_1_weights[5][0] = 11;
        layer_1_weights[6][0] = 0;
        layer_1_weights[7][0] = 1;
        layer_1_weights[8][0] = 3;
        layer_1_weights[9][0] = 36;
        layer_1_weights[10][0] = -1;
        layer_1_weights[11][0] = 1;
        layer_1_weights[12][0] = 2;
        layer_1_weights[13][0] = -2;
        layer_1_weights[14][0] = -10;
        layer_1_weights[15][0] = 1;
        layer_1_weights[16][0] = 6;
        layer_1_weights[17][0] = 2;
        layer_1_weights[18][0] = 3;
        layer_1_weights[19][0] = 3;
        layer_1_weights[20][0] = 6;
        layer_1_weights[21][0] = 7;
        layer_1_weights[22][0] = 16;
        layer_1_weights[23][0] = 9;
        layer_1_weights[24][0] = 2;
        layer_1_weights[25][0] = -10;
        layer_1_weights[26][0] = -2;
        layer_1_weights[27][0] = 1;
        layer_1_weights[28][0] = -2;
        layer_1_weights[29][0] = -2;
        layer_1_weights[30][0] = 1;
        layer_1_weights[31][0] = 1;
        layer_1_weights[32][0] = 3;
        layer_1_weights[33][0] = 4;
        layer_1_weights[34][0] = 10;
        layer_1_weights[35][0] = 38;
        layer_1_weights[36][0] = -16;
        layer_1_weights[37][0] = -4;
        layer_1_weights[38][0] = -6;
        layer_1_weights[39][0] = 1;
        layer_1_weights[40][0] = -1;
        layer_1_weights[41][0] = 1;
        layer_1_weights[42][0] = -6;
        layer_1_weights[43][0] = -4;
        layer_1_weights[44][0] = 2;
        layer_1_weights[45][0] = 4;
        layer_1_weights[46][0] = 12;
        layer_1_weights[47][0] = 39;
        layer_1_weights[48][0] = -31;
        layer_1_weights[49][0] = 0;
        layer_1_weights[50][0] = -4;
        layer_1_weights[51][0] = 6;
        layer_1_weights[52][0] = 9;
        layer_1_weights[53][0] = 12;
        layer_1_weights[54][0] = -6;
        layer_1_weights[55][0] = -7;
        layer_1_weights[56][0] = 1;
        layer_1_weights[57][0] = 6;
        layer_1_weights[58][0] = 16;
        layer_1_weights[59][0] = 16;
        layer_1_weights[60][0] = -29;
        layer_1_weights[61][0] = -7;
        layer_1_weights[62][0] = 13;
        layer_1_weights[63][0] = 10;
        layer_1_weights[64][0] = 9;
        layer_1_weights[65][0] = 13;
        layer_1_weights[66][0] = 5;
        layer_1_weights[67][0] = 0;
        layer_1_weights[68][0] = 2;
        layer_1_weights[69][0] = 10;
        layer_1_weights[70][0] = 11;
        layer_1_weights[71][0] = -17;
        layer_1_weights[72][0] = -7;
        layer_1_weights[73][0] = -11;
        layer_1_weights[74][0] = -4;
        layer_1_weights[75][0] = -3;
        layer_1_weights[76][0] = 2;
        layer_1_weights[77][0] = 11;
        layer_1_weights[78][0] = 0;
        layer_1_weights[79][0] = -5;
        layer_1_weights[80][0] = -5;
        layer_1_weights[81][0] = 0;
        layer_1_weights[82][0] = 2;
        layer_1_weights[83][0] = -14;
        layer_1_weights[84][0] = -9;
        layer_1_weights[85][0] = -13;
        layer_1_weights[86][0] = -4;
        layer_1_weights[87][0] = 0;
        layer_1_weights[88][0] = 11;
        layer_1_weights[89][0] = 2;
        layer_1_weights[90][0] = -8;
        layer_1_weights[91][0] = -4;
        layer_1_weights[92][0] = -6;
        layer_1_weights[93][0] = -2;
        layer_1_weights[94][0] = -5;
        layer_1_weights[95][0] = -20;
        layer_1_weights[96][0] = 9;
        layer_1_weights[97][0] = -7;
        layer_1_weights[98][0] = -1;
        layer_1_weights[99][0] = 4;
        layer_1_weights[100][0] = 9;
        layer_1_weights[101][0] = 2;
        layer_1_weights[102][0] = -2;
        layer_1_weights[103][0] = 2;
        layer_1_weights[104][0] = 1;
        layer_1_weights[105][0] = -2;
        layer_1_weights[106][0] = -3;
        layer_1_weights[107][0] = -24;
        layer_1_weights[108][0] = -14;
        layer_1_weights[109][0] = -13;
        layer_1_weights[110][0] = -3;
        layer_1_weights[111][0] = -1;
        layer_1_weights[112][0] = 1;
        layer_1_weights[113][0] = 17;
        layer_1_weights[114][0] = 14;
        layer_1_weights[115][0] = 4;
        layer_1_weights[116][0] = -2;
        layer_1_weights[117][0] = -3;
        layer_1_weights[118][0] = -5;
        layer_1_weights[119][0] = 8;
        layer_1_weights[120][0] = -3;
        layer_1_weights[121][0] = -15;
        layer_1_weights[122][0] = -8;
        layer_1_weights[123][0] = -1;
        layer_1_weights[124][0] = -1;
        layer_1_weights[125][0] = 8;
        layer_1_weights[126][0] = 7;
        layer_1_weights[127][0] = 3;
        layer_1_weights[128][0] = -2;
        layer_1_weights[129][0] = -2;
        layer_1_weights[130][0] = -8;
        layer_1_weights[131][0] = -15;
        layer_1_weights[132][0] = -1;
        layer_1_weights[133][0] = -3;
        layer_1_weights[134][0] = -6;
        layer_1_weights[135][0] = -12;
        layer_1_weights[136][0] = -6;
        layer_1_weights[137][0] = -3;
        layer_1_weights[138][0] = -1;
        layer_1_weights[139][0] = -1;
        layer_1_weights[140][0] = 4;
        layer_1_weights[141][0] = -4;
        layer_1_weights[142][0] = -2;
        layer_1_weights[143][0] = -3;
        layer_1_weights[0][1] = 1;
        layer_1_weights[1][1] = -3;
        layer_1_weights[2][1] = -18;
        layer_1_weights[3][1] = -18;
        layer_1_weights[4][1] = -14;
        layer_1_weights[5][1] = -16;
        layer_1_weights[6][1] = 4;
        layer_1_weights[7][1] = -7;
        layer_1_weights[8][1] = 3;
        layer_1_weights[9][1] = -25;
        layer_1_weights[10][1] = 2;
        layer_1_weights[11][1] = 1;
        layer_1_weights[12][1] = 1;
        layer_1_weights[13][1] = 1;
        layer_1_weights[14][1] = -2;
        layer_1_weights[15][1] = -2;
        layer_1_weights[16][1] = -2;
        layer_1_weights[17][1] = -6;
        layer_1_weights[18][1] = -6;
        layer_1_weights[19][1] = -2;
        layer_1_weights[20][1] = -5;
        layer_1_weights[21][1] = -7;
        layer_1_weights[22][1] = -7;
        layer_1_weights[23][1] = 3;
        layer_1_weights[24][1] = -3;
        layer_1_weights[25][1] = 7;
        layer_1_weights[26][1] = 12;
        layer_1_weights[27][1] = 9;
        layer_1_weights[28][1] = 8;
        layer_1_weights[29][1] = 8;
        layer_1_weights[30][1] = 4;
        layer_1_weights[31][1] = 1;
        layer_1_weights[32][1] = 1;
        layer_1_weights[33][1] = -1;
        layer_1_weights[34][1] = -3;
        layer_1_weights[35][1] = 7;
        layer_1_weights[36][1] = 16;
        layer_1_weights[37][1] = 14;
        layer_1_weights[38][1] = 15;
        layer_1_weights[39][1] = 10;
        layer_1_weights[40][1] = 6;
        layer_1_weights[41][1] = 3;
        layer_1_weights[42][1] = 3;
        layer_1_weights[43][1] = 10;
        layer_1_weights[44][1] = 7;
        layer_1_weights[45][1] = 5;
        layer_1_weights[46][1] = 4;
        layer_1_weights[47][1] = 2;
        layer_1_weights[48][1] = 12;
        layer_1_weights[49][1] = 21;
        layer_1_weights[50][1] = 6;
        layer_1_weights[51][1] = 1;
        layer_1_weights[52][1] = -1;
        layer_1_weights[53][1] = 7;
        layer_1_weights[54][1] = 2;
        layer_1_weights[55][1] = 11;
        layer_1_weights[56][1] = 11;
        layer_1_weights[57][1] = 10;
        layer_1_weights[58][1] = 12;
        layer_1_weights[59][1] = 15;
        layer_1_weights[60][1] = 12;
        layer_1_weights[61][1] = 0;
        layer_1_weights[62][1] = -8;
        layer_1_weights[63][1] = 0;
        layer_1_weights[64][1] = 6;
        layer_1_weights[65][1] = 4;
        layer_1_weights[66][1] = 0;
        layer_1_weights[67][1] = 5;
        layer_1_weights[68][1] = 3;
        layer_1_weights[69][1] = 2;
        layer_1_weights[70][1] = -10;
        layer_1_weights[71][1] = 11;
        layer_1_weights[72][1] = -3;
        layer_1_weights[73][1] = 14;
        layer_1_weights[74][1] = 3;
        layer_1_weights[75][1] = 4;
        layer_1_weights[76][1] = -1;
        layer_1_weights[77][1] = -2;
        layer_1_weights[78][1] = -12;
        layer_1_weights[79][1] = 2;
        layer_1_weights[80][1] = 9;
        layer_1_weights[81][1] = 2;
        layer_1_weights[82][1] = 5;
        layer_1_weights[83][1] = 3;
        layer_1_weights[84][1] = 23;
        layer_1_weights[85][1] = 15;
        layer_1_weights[86][1] = 7;
        layer_1_weights[87][1] = -1;
        layer_1_weights[88][1] = -5;
        layer_1_weights[89][1] = -8;
        layer_1_weights[90][1] = -3;
        layer_1_weights[91][1] = 5;
        layer_1_weights[92][1] = 2;
        layer_1_weights[93][1] = -2;
        layer_1_weights[94][1] = 0;
        layer_1_weights[95][1] = -5;
        layer_1_weights[96][1] = 17;
        layer_1_weights[97][1] = 19;
        layer_1_weights[98][1] = 3;
        layer_1_weights[99][1] = -2;
        layer_1_weights[100][1] = -8;
        layer_1_weights[101][1] = -11;
        layer_1_weights[102][1] = -4;
        layer_1_weights[103][1] = -2;
        layer_1_weights[104][1] = -4;
        layer_1_weights[105][1] = -5;
        layer_1_weights[106][1] = -9;
        layer_1_weights[107][1] = -14;
        layer_1_weights[108][1] = 7;
        layer_1_weights[109][1] = -8;
        layer_1_weights[110][1] = 0;
        layer_1_weights[111][1] = -2;
        layer_1_weights[112][1] = 1;
        layer_1_weights[113][1] = 3;
        layer_1_weights[114][1] = 3;
        layer_1_weights[115][1] = -2;
        layer_1_weights[116][1] = -5;
        layer_1_weights[117][1] = -11;
        layer_1_weights[118][1] = -12;
        layer_1_weights[119][1] = -16;
        layer_1_weights[120][1] = 0;
        layer_1_weights[121][1] = 16;
        layer_1_weights[122][1] = 4;
        layer_1_weights[123][1] = 6;
        layer_1_weights[124][1] = 6;
        layer_1_weights[125][1] = 8;
        layer_1_weights[126][1] = 5;
        layer_1_weights[127][1] = 1;
        layer_1_weights[128][1] = -2;
        layer_1_weights[129][1] = -6;
        layer_1_weights[130][1] = -7;
        layer_1_weights[131][1] = 0;
        layer_1_weights[132][1] = -2;
        layer_1_weights[133][1] = 6;
        layer_1_weights[134][1] = 5;
        layer_1_weights[135][1] = 20;
        layer_1_weights[136][1] = 23;
        layer_1_weights[137][1] = 23;
        layer_1_weights[138][1] = 22;
        layer_1_weights[139][1] = 21;
        layer_1_weights[140][1] = 16;
        layer_1_weights[141][1] = 11;
        layer_1_weights[142][1] = -3;
        layer_1_weights[143][1] = 1;
        layer_1_weights[0][2] = 1;
        layer_1_weights[1][2] = -1;
        layer_1_weights[2][2] = 1;
        layer_1_weights[3][2] = 4;
        layer_1_weights[4][2] = -15;
        layer_1_weights[5][2] = 0;
        layer_1_weights[6][2] = 6;
        layer_1_weights[7][2] = 7;
        layer_1_weights[8][2] = -2;
        layer_1_weights[9][2] = -13;
        layer_1_weights[10][2] = 2;
        layer_1_weights[11][2] = 0;
        layer_1_weights[12][2] = -3;
        layer_1_weights[13][2] = 1;
        layer_1_weights[14][2] = 18;
        layer_1_weights[15][2] = 13;
        layer_1_weights[16][2] = 15;
        layer_1_weights[17][2] = 11;
        layer_1_weights[18][2] = 10;
        layer_1_weights[19][2] = 6;
        layer_1_weights[20][2] = 0;
        layer_1_weights[21][2] = -3;
        layer_1_weights[22][2] = -9;
        layer_1_weights[23][2] = -3;
        layer_1_weights[24][2] = -3;
        layer_1_weights[25][2] = 6;
        layer_1_weights[26][2] = 4;
        layer_1_weights[27][2] = 3;
        layer_1_weights[28][2] = 4;
        layer_1_weights[29][2] = 7;
        layer_1_weights[30][2] = 3;
        layer_1_weights[31][2] = 0;
        layer_1_weights[32][2] = 0;
        layer_1_weights[33][2] = -2;
        layer_1_weights[34][2] = -2;
        layer_1_weights[35][2] = 11;
        layer_1_weights[36][2] = -7;
        layer_1_weights[37][2] = 7;
        layer_1_weights[38][2] = 4;
        layer_1_weights[39][2] = 2;
        layer_1_weights[40][2] = -2;
        layer_1_weights[41][2] = -3;
        layer_1_weights[42][2] = 1;
        layer_1_weights[43][2] = 0;
        layer_1_weights[44][2] = -1;
        layer_1_weights[45][2] = 0;
        layer_1_weights[46][2] = 0;
        layer_1_weights[47][2] = 9;
        layer_1_weights[48][2] = 8;
        layer_1_weights[49][2] = 5;
        layer_1_weights[50][2] = 0;
        layer_1_weights[51][2] = -2;
        layer_1_weights[52][2] = -7;
        layer_1_weights[53][2] = 0;
        layer_1_weights[54][2] = 6;
        layer_1_weights[55][2] = -1;
        layer_1_weights[56][2] = 2;
        layer_1_weights[57][2] = -2;
        layer_1_weights[58][2] = 9;
        layer_1_weights[59][2] = 12;
        layer_1_weights[60][2] = -32;
        layer_1_weights[61][2] = 5;
        layer_1_weights[62][2] = -6;
        layer_1_weights[63][2] = -3;
        layer_1_weights[64][2] = -3;
        layer_1_weights[65][2] = 15;
        layer_1_weights[66][2] = 20;
        layer_1_weights[67][2] = 3;
        layer_1_weights[68][2] = -1;
        layer_1_weights[69][2] = -9;
        layer_1_weights[70][2] = -5;
        layer_1_weights[71][2] = -4;
        layer_1_weights[72][2] = 6;
        layer_1_weights[73][2] = -10;
        layer_1_weights[74][2] = -6;
        layer_1_weights[75][2] = -8;
        layer_1_weights[76][2] = -1;
        layer_1_weights[77][2] = 11;
        layer_1_weights[78][2] = 12;
        layer_1_weights[79][2] = -3;
        layer_1_weights[80][2] = -6;
        layer_1_weights[81][2] = -5;
        layer_1_weights[82][2] = -4;
        layer_1_weights[83][2] = -8;
        layer_1_weights[84][2] = 24;
        layer_1_weights[85][2] = 2;
        layer_1_weights[86][2] = -5;
        layer_1_weights[87][2] = -12;
        layer_1_weights[88][2] = -9;
        layer_1_weights[89][2] = -7;
        layer_1_weights[90][2] = -5;
        layer_1_weights[91][2] = -4;
        layer_1_weights[92][2] = 0;
        layer_1_weights[93][2] = 1;
        layer_1_weights[94][2] = -5;
        layer_1_weights[95][2] = 12;
        layer_1_weights[96][2] = -3;
        layer_1_weights[97][2] = 3;
        layer_1_weights[98][2] = 10;
        layer_1_weights[99][2] = 7;
        layer_1_weights[100][2] = -4;
        layer_1_weights[101][2] = -4;
        layer_1_weights[102][2] = -3;
        layer_1_weights[103][2] = 4;
        layer_1_weights[104][2] = 5;
        layer_1_weights[105][2] = 4;
        layer_1_weights[106][2] = 3;
        layer_1_weights[107][2] = 1;
        layer_1_weights[108][2] = 15;
        layer_1_weights[109][2] = 6;
        layer_1_weights[110][2] = 7;
        layer_1_weights[111][2] = 7;
        layer_1_weights[112][2] = 2;
        layer_1_weights[113][2] = 1;
        layer_1_weights[114][2] = 5;
        layer_1_weights[115][2] = 5;
        layer_1_weights[116][2] = 4;
        layer_1_weights[117][2] = 1;
        layer_1_weights[118][2] = -9;
        layer_1_weights[119][2] = -8;
        layer_1_weights[120][2] = -2;
        layer_1_weights[121][2] = 5;
        layer_1_weights[122][2] = 3;
        layer_1_weights[123][2] = 2;
        layer_1_weights[124][2] = 3;
        layer_1_weights[125][2] = 5;
        layer_1_weights[126][2] = 2;
        layer_1_weights[127][2] = 0;
        layer_1_weights[128][2] = 0;
        layer_1_weights[129][2] = -7;
        layer_1_weights[130][2] = -5;
        layer_1_weights[131][2] = -12;
        layer_1_weights[132][2] = 1;
        layer_1_weights[133][2] = -2;
        layer_1_weights[134][2] = 8;
        layer_1_weights[135][2] = 16;
        layer_1_weights[136][2] = 13;
        layer_1_weights[137][2] = 5;
        layer_1_weights[138][2] = 7;
        layer_1_weights[139][2] = 7;
        layer_1_weights[140][2] = 0;
        layer_1_weights[141][2] = 20;
        layer_1_weights[142][2] = 0;
        layer_1_weights[143][2] = 2;
        layer_1_weights[0][3] = 0;
        layer_1_weights[1][3] = 3;
        layer_1_weights[2][3] = 20;
        layer_1_weights[3][3] = 9;
        layer_1_weights[4][3] = 4;
        layer_1_weights[5][3] = 3;
        layer_1_weights[6][3] = 5;
        layer_1_weights[7][3] = -10;
        layer_1_weights[8][3] = 7;
        layer_1_weights[9][3] = 8;
        layer_1_weights[10][3] = 0;
        layer_1_weights[11][3] = -2;
        layer_1_weights[12][3] = 3;
        layer_1_weights[13][3] = 3;
        layer_1_weights[14][3] = 22;
        layer_1_weights[15][3] = 5;
        layer_1_weights[16][3] = -1;
        layer_1_weights[17][3] = 1;
        layer_1_weights[18][3] = 1;
        layer_1_weights[19][3] = -3;
        layer_1_weights[20][3] = -1;
        layer_1_weights[21][3] = -2;
        layer_1_weights[22][3] = -5;
        layer_1_weights[23][3] = -9;
        layer_1_weights[24][3] = 0;
        layer_1_weights[25][3] = 21;
        layer_1_weights[26][3] = 6;
        layer_1_weights[27][3] = 4;
        layer_1_weights[28][3] = 0;
        layer_1_weights[29][3] = 1;
        layer_1_weights[30][3] = 1;
        layer_1_weights[31][3] = -2;
        layer_1_weights[32][3] = -3;
        layer_1_weights[33][3] = -3;
        layer_1_weights[34][3] = -2;
        layer_1_weights[35][3] = 2;
        layer_1_weights[36][3] = 10;
        layer_1_weights[37][3] = 14;
        layer_1_weights[38][3] = 5;
        layer_1_weights[39][3] = 2;
        layer_1_weights[40][3] = -2;
        layer_1_weights[41][3] = 1;
        layer_1_weights[42][3] = 3;
        layer_1_weights[43][3] = 2;
        layer_1_weights[44][3] = -4;
        layer_1_weights[45][3] = -4;
        layer_1_weights[46][3] = -17;
        layer_1_weights[47][3] = 2;
        layer_1_weights[48][3] = 15;
        layer_1_weights[49][3] = 1;
        layer_1_weights[50][3] = -3;
        layer_1_weights[51][3] = -1;
        layer_1_weights[52][3] = -2;
        layer_1_weights[53][3] = 2;
        layer_1_weights[54][3] = 8;
        layer_1_weights[55][3] = 6;
        layer_1_weights[56][3] = 8;
        layer_1_weights[57][3] = 3;
        layer_1_weights[58][3] = -18;
        layer_1_weights[59][3] = -20;
        layer_1_weights[60][3] = 10;
        layer_1_weights[61][3] = 7;
        layer_1_weights[62][3] = 4;
        layer_1_weights[63][3] = 3;
        layer_1_weights[64][3] = -2;
        layer_1_weights[65][3] = -1;
        layer_1_weights[66][3] = 15;
        layer_1_weights[67][3] = 14;
        layer_1_weights[68][3] = 10;
        layer_1_weights[69][3] = 21;
        layer_1_weights[70][3] = -1;
        layer_1_weights[71][3] = -48;
        layer_1_weights[72][3] = -3;
        layer_1_weights[73][3] = -2;
        layer_1_weights[74][3] = 2;
        layer_1_weights[75][3] = -5;
        layer_1_weights[76][3] = -2;
        layer_1_weights[77][3] = 5;
        layer_1_weights[78][3] = 16;
        layer_1_weights[79][3] = 8;
        layer_1_weights[80][3] = 0;
        layer_1_weights[81][3] = 0;
        layer_1_weights[82][3] = -5;
        layer_1_weights[83][3] = -3;
        layer_1_weights[84][3] = 23;
        layer_1_weights[85][3] = -18;
        layer_1_weights[86][3] = -13;
        layer_1_weights[87][3] = 2;
        layer_1_weights[88][3] = 7;
        layer_1_weights[89][3] = 4;
        layer_1_weights[90][3] = 6;
        layer_1_weights[91][3] = -4;
        layer_1_weights[92][3] = -3;
        layer_1_weights[93][3] = -6;
        layer_1_weights[94][3] = -14;
        layer_1_weights[95][3] = -4;
        layer_1_weights[96][3] = -12;
        layer_1_weights[97][3] = -12;
        layer_1_weights[98][3] = -9;
        layer_1_weights[99][3] = -7;
        layer_1_weights[100][3] = 0;
        layer_1_weights[101][3] = -1;
        layer_1_weights[102][3] = -4;
        layer_1_weights[103][3] = -4;
        layer_1_weights[104][3] = -4;
        layer_1_weights[105][3] = -8;
        layer_1_weights[106][3] = -17;
        layer_1_weights[107][3] = 9;
        layer_1_weights[108][3] = 5;
        layer_1_weights[109][3] = -6;
        layer_1_weights[110][3] = -2;
        layer_1_weights[111][3] = -5;
        layer_1_weights[112][3] = -7;
        layer_1_weights[113][3] = 3;
        layer_1_weights[114][3] = 3;
        layer_1_weights[115][3] = 0;
        layer_1_weights[116][3] = -7;
        layer_1_weights[117][3] = -10;
        layer_1_weights[118][3] = -16;
        layer_1_weights[119][3] = -4;
        layer_1_weights[120][3] = 3;
        layer_1_weights[121][3] = -12;
        layer_1_weights[122][3] = 3;
        layer_1_weights[123][3] = 2;
        layer_1_weights[124][3] = -2;
        layer_1_weights[125][3] = 1;
        layer_1_weights[126][3] = 0;
        layer_1_weights[127][3] = -3;
        layer_1_weights[128][3] = -4;
        layer_1_weights[129][3] = -7;
        layer_1_weights[130][3] = -3;
        layer_1_weights[131][3] = -17;
        layer_1_weights[132][3] = -1;
        layer_1_weights[133][3] = 24;
        layer_1_weights[134][3] = 9;
        layer_1_weights[135][3] = 7;
        layer_1_weights[136][3] = 0;
        layer_1_weights[137][3] = -5;
        layer_1_weights[138][3] = 2;
        layer_1_weights[139][3] = 3;
        layer_1_weights[140][3] = 6;
        layer_1_weights[141][3] = 9;
        layer_1_weights[142][3] = 1;
        layer_1_weights[143][3] = -2;
        layer_1_weights[0][4] = -2;
        layer_1_weights[1][4] = 0;
        layer_1_weights[2][4] = -17;
        layer_1_weights[3][4] = -15;
        layer_1_weights[4][4] = -10;
        layer_1_weights[5][4] = -14;
        layer_1_weights[6][4] = -12;
        layer_1_weights[7][4] = -9;
        layer_1_weights[8][4] = -11;
        layer_1_weights[9][4] = -25;
        layer_1_weights[10][4] = -3;
        layer_1_weights[11][4] = -2;
        layer_1_weights[12][4] = -3;
        layer_1_weights[13][4] = 3;
        layer_1_weights[14][4] = 0;
        layer_1_weights[15][4] = 5;
        layer_1_weights[16][4] = 7;
        layer_1_weights[17][4] = 6;
        layer_1_weights[18][4] = 4;
        layer_1_weights[19][4] = 1;
        layer_1_weights[20][4] = 1;
        layer_1_weights[21][4] = 0;
        layer_1_weights[22][4] = 3;
        layer_1_weights[23][4] = -8;
        layer_1_weights[24][4] = -2;
        layer_1_weights[25][4] = 6;
        layer_1_weights[26][4] = 1;
        layer_1_weights[27][4] = 3;
        layer_1_weights[28][4] = 0;
        layer_1_weights[29][4] = 2;
        layer_1_weights[30][4] = 6;
        layer_1_weights[31][4] = 3;
        layer_1_weights[32][4] = 0;
        layer_1_weights[33][4] = 2;
        layer_1_weights[34][4] = 3;
        layer_1_weights[35][4] = -6;
        layer_1_weights[36][4] = -8;
        layer_1_weights[37][4] = 5;
        layer_1_weights[38][4] = 0;
        layer_1_weights[39][4] = -2;
        layer_1_weights[40][4] = 0;
        layer_1_weights[41][4] = 0;
        layer_1_weights[42][4] = -4;
        layer_1_weights[43][4] = 0;
        layer_1_weights[44][4] = 1;
        layer_1_weights[45][4] = -2;
        layer_1_weights[46][4] = -3;
        layer_1_weights[47][4] = 6;
        layer_1_weights[48][4] = -17;
        layer_1_weights[49][4] = -2;
        layer_1_weights[50][4] = 2;
        layer_1_weights[51][4] = -1;
        layer_1_weights[52][4] = 3;
        layer_1_weights[53][4] = -5;
        layer_1_weights[54][4] = -10;
        layer_1_weights[55][4] = 0;
        layer_1_weights[56][4] = 4;
        layer_1_weights[57][4] = 3;
        layer_1_weights[58][4] = -2;
        layer_1_weights[59][4] = -11;
        layer_1_weights[60][4] = -3;
        layer_1_weights[61][4] = 0;
        layer_1_weights[62][4] = -4;
        layer_1_weights[63][4] = 0;
        layer_1_weights[64][4] = 6;
        layer_1_weights[65][4] = 0;
        layer_1_weights[66][4] = -4;
        layer_1_weights[67][4] = 9;
        layer_1_weights[68][4] = 6;
        layer_1_weights[69][4] = 10;
        layer_1_weights[70][4] = 4;
        layer_1_weights[71][4] = 8;
        layer_1_weights[72][4] = 5;
        layer_1_weights[73][4] = -1;
        layer_1_weights[74][4] = 1;
        layer_1_weights[75][4] = 8;
        layer_1_weights[76][4] = 5;
        layer_1_weights[77][4] = 17;
        layer_1_weights[78][4] = 7;
        layer_1_weights[79][4] = 8;
        layer_1_weights[80][4] = 2;
        layer_1_weights[81][4] = -3;
        layer_1_weights[82][4] = 1;
        layer_1_weights[83][4] = 19;
        layer_1_weights[84][4] = -17;
        layer_1_weights[85][4] = 5;
        layer_1_weights[86][4] = 7;
        layer_1_weights[87][4] = 7;
        layer_1_weights[88][4] = 7;
        layer_1_weights[89][4] = 11;
        layer_1_weights[90][4] = 8;
        layer_1_weights[91][4] = 3;
        layer_1_weights[92][4] = -3;
        layer_1_weights[93][4] = -3;
        layer_1_weights[94][4] = 4;
        layer_1_weights[95][4] = 4;
        layer_1_weights[96][4] = -10;
        layer_1_weights[97][4] = 5;
        layer_1_weights[98][4] = 4;
        layer_1_weights[99][4] = -2;
        layer_1_weights[100][4] = 0;
        layer_1_weights[101][4] = -4;
        layer_1_weights[102][4] = 0;
        layer_1_weights[103][4] = 2;
        layer_1_weights[104][4] = 1;
        layer_1_weights[105][4] = 2;
        layer_1_weights[106][4] = -1;
        layer_1_weights[107][4] = 7;
        layer_1_weights[108][4] = 17;
        layer_1_weights[109][4] = -7;
        layer_1_weights[110][4] = -7;
        layer_1_weights[111][4] = -3;
        layer_1_weights[112][4] = -2;
        layer_1_weights[113][4] = 1;
        layer_1_weights[114][4] = 0;
        layer_1_weights[115][4] = 0;
        layer_1_weights[116][4] = 4;
        layer_1_weights[117][4] = 1;
        layer_1_weights[118][4] = 0;
        layer_1_weights[119][4] = -11;
        layer_1_weights[120][4] = -2;
        layer_1_weights[121][4] = -4;
        layer_1_weights[122][4] = -9;
        layer_1_weights[123][4] = -4;
        layer_1_weights[124][4] = -4;
        layer_1_weights[125][4] = -3;
        layer_1_weights[126][4] = -5;
        layer_1_weights[127][4] = 2;
        layer_1_weights[128][4] = 7;
        layer_1_weights[129][4] = 16;
        layer_1_weights[130][4] = 9;
        layer_1_weights[131][4] = 12;
        layer_1_weights[132][4] = 2;
        layer_1_weights[133][4] = -2;
        layer_1_weights[134][4] = 0;
        layer_1_weights[135][4] = -4;
        layer_1_weights[136][4] = -2;
        layer_1_weights[137][4] = 0;
        layer_1_weights[138][4] = -2;
        layer_1_weights[139][4] = 0;
        layer_1_weights[140][4] = -6;
        layer_1_weights[141][4] = -8;
        layer_1_weights[142][4] = -1;
        layer_1_weights[143][4] = -2;
        layer_1_weights[0][5] = -2;
        layer_1_weights[1][5] = 1;
        layer_1_weights[2][5] = 14;
        layer_1_weights[3][5] = 29;
        layer_1_weights[4][5] = 31;
        layer_1_weights[5][5] = 24;
        layer_1_weights[6][5] = 5;
        layer_1_weights[7][5] = 33;
        layer_1_weights[8][5] = 5;
        layer_1_weights[9][5] = 39;
        layer_1_weights[10][5] = 1;
        layer_1_weights[11][5] = 2;
        layer_1_weights[12][5] = 2;
        layer_1_weights[13][5] = -2;
        layer_1_weights[14][5] = 19;
        layer_1_weights[15][5] = 18;
        layer_1_weights[16][5] = 27;
        layer_1_weights[17][5] = 14;
        layer_1_weights[18][5] = 12;
        layer_1_weights[19][5] = 13;
        layer_1_weights[20][5] = 7;
        layer_1_weights[21][5] = -1;
        layer_1_weights[22][5] = -7;
        layer_1_weights[23][5] = 1;
        layer_1_weights[24][5] = -2;
        layer_1_weights[25][5] = 6;
        layer_1_weights[26][5] = 17;
        layer_1_weights[27][5] = 12;
        layer_1_weights[28][5] = 3;
        layer_1_weights[29][5] = 3;
        layer_1_weights[30][5] = 2;
        layer_1_weights[31][5] = -3;
        layer_1_weights[32][5] = -3;
        layer_1_weights[33][5] = -3;
        layer_1_weights[34][5] = -2;
        layer_1_weights[35][5] = 5;
        layer_1_weights[36][5] = 10;
        layer_1_weights[37][5] = 25;
        layer_1_weights[38][5] = 2;
        layer_1_weights[39][5] = 2;
        layer_1_weights[40][5] = -3;
        layer_1_weights[41][5] = -8;
        layer_1_weights[42][5] = -3;
        layer_1_weights[43][5] = -5;
        layer_1_weights[44][5] = -4;
        layer_1_weights[45][5] = -6;
        layer_1_weights[46][5] = -7;
        layer_1_weights[47][5] = -5;
        layer_1_weights[48][5] = 15;
        layer_1_weights[49][5] = 12;
        layer_1_weights[50][5] = -9;
        layer_1_weights[51][5] = -11;
        layer_1_weights[52][5] = -12;
        layer_1_weights[53][5] = -4;
        layer_1_weights[54][5] = 0;
        layer_1_weights[55][5] = -3;
        layer_1_weights[56][5] = 0;
        layer_1_weights[57][5] = 2;
        layer_1_weights[58][5] = -3;
        layer_1_weights[59][5] = -12;
        layer_1_weights[60][5] = -11;
        layer_1_weights[61][5] = -15;
        layer_1_weights[62][5] = -13;
        layer_1_weights[63][5] = -9;
        layer_1_weights[64][5] = -1;
        layer_1_weights[65][5] = 7;
        layer_1_weights[66][5] = 5;
        layer_1_weights[67][5] = -5;
        layer_1_weights[68][5] = 1;
        layer_1_weights[69][5] = 7;
        layer_1_weights[70][5] = 9;
        layer_1_weights[71][5] = 7;
        layer_1_weights[72][5] = -12;
        layer_1_weights[73][5] = -6;
        layer_1_weights[74][5] = 5;
        layer_1_weights[75][5] = 8;
        layer_1_weights[76][5] = 13;
        layer_1_weights[77][5] = 8;
        layer_1_weights[78][5] = 2;
        layer_1_weights[79][5] = -2;
        layer_1_weights[80][5] = 2;
        layer_1_weights[81][5] = 5;
        layer_1_weights[82][5] = 12;
        layer_1_weights[83][5] = 28;
        layer_1_weights[84][5] = 14;
        layer_1_weights[85][5] = 11;
        layer_1_weights[86][5] = 5;
        layer_1_weights[87][5] = 2;
        layer_1_weights[88][5] = 4;
        layer_1_weights[89][5] = -1;
        layer_1_weights[90][5] = -3;
        layer_1_weights[91][5] = 4;
        layer_1_weights[92][5] = 8;
        layer_1_weights[93][5] = 4;
        layer_1_weights[94][5] = 10;
        layer_1_weights[95][5] = 17;
        layer_1_weights[96][5] = 16;
        layer_1_weights[97][5] = 8;
        layer_1_weights[98][5] = 7;
        layer_1_weights[99][5] = 3;
        layer_1_weights[100][5] = 9;
        layer_1_weights[101][5] = 2;
        layer_1_weights[102][5] = 6;
        layer_1_weights[103][5] = 12;
        layer_1_weights[104][5] = 8;
        layer_1_weights[105][5] = 9;
        layer_1_weights[106][5] = -2;
        layer_1_weights[107][5] = 9;
        layer_1_weights[108][5] = 15;
        layer_1_weights[109][5] = -2;
        layer_1_weights[110][5] = -3;
        layer_1_weights[111][5] = 3;
        layer_1_weights[112][5] = 6;
        layer_1_weights[113][5] = 9;
        layer_1_weights[114][5] = 9;
        layer_1_weights[115][5] = 4;
        layer_1_weights[116][5] = 1;
        layer_1_weights[117][5] = -7;
        layer_1_weights[118][5] = -10;
        layer_1_weights[119][5] = -2;
        layer_1_weights[120][5] = 2;
        layer_1_weights[121][5] = 7;
        layer_1_weights[122][5] = 1;
        layer_1_weights[123][5] = 1;
        layer_1_weights[124][5] = -3;
        layer_1_weights[125][5] = 0;
        layer_1_weights[126][5] = -4;
        layer_1_weights[127][5] = -8;
        layer_1_weights[128][5] = -12;
        layer_1_weights[129][5] = -12;
        layer_1_weights[130][5] = -18;
        layer_1_weights[131][5] = 3;
        layer_1_weights[132][5] = 2;
        layer_1_weights[133][5] = -7;
        layer_1_weights[134][5] = -25;
        layer_1_weights[135][5] = -13;
        layer_1_weights[136][5] = -10;
        layer_1_weights[137][5] = -13;
        layer_1_weights[138][5] = -13;
        layer_1_weights[139][5] = -12;
        layer_1_weights[140][5] = -22;
        layer_1_weights[141][5] = -24;
        layer_1_weights[142][5] = 0;
        layer_1_weights[143][5] = -2;
        layer_1_weights[0][6] = 0;
        layer_1_weights[1][6] = 3;
        layer_1_weights[2][6] = 0;
        layer_1_weights[3][6] = 9;
        layer_1_weights[4][6] = 12;
        layer_1_weights[5][6] = 21;
        layer_1_weights[6][6] = 10;
        layer_1_weights[7][6] = -2;
        layer_1_weights[8][6] = 0;
        layer_1_weights[9][6] = 3;
        layer_1_weights[10][6] = 2;
        layer_1_weights[11][6] = -2;
        layer_1_weights[12][6] = 1;
        layer_1_weights[13][6] = 0;
        layer_1_weights[14][6] = 4;
        layer_1_weights[15][6] = 10;
        layer_1_weights[16][6] = 5;
        layer_1_weights[17][6] = 10;
        layer_1_weights[18][6] = 6;
        layer_1_weights[19][6] = -2;
        layer_1_weights[20][6] = -5;
        layer_1_weights[21][6] = -3;
        layer_1_weights[22][6] = -17;
        layer_1_weights[23][6] = -8;
        layer_1_weights[24][6] = -1;
        layer_1_weights[25][6] = 8;
        layer_1_weights[26][6] = -14;
        layer_1_weights[27][6] = -2;
        layer_1_weights[28][6] = 0;
        layer_1_weights[29][6] = 4;
        layer_1_weights[30][6] = 8;
        layer_1_weights[31][6] = 4;
        layer_1_weights[32][6] = 1;
        layer_1_weights[33][6] = -4;
        layer_1_weights[34][6] = -10;
        layer_1_weights[35][6] = -7;
        layer_1_weights[36][6] = 3;
        layer_1_weights[37][6] = -5;
        layer_1_weights[38][6] = -3;
        layer_1_weights[39][6] = 0;
        layer_1_weights[40][6] = 2;
        layer_1_weights[41][6] = 12;
        layer_1_weights[42][6] = 18;
        layer_1_weights[43][6] = 14;
        layer_1_weights[44][6] = 2;
        layer_1_weights[45][6] = -2;
        layer_1_weights[46][6] = -5;
        layer_1_weights[47][6] = -19;
        layer_1_weights[48][6] = -18;
        layer_1_weights[49][6] = 1;
        layer_1_weights[50][6] = 3;
        layer_1_weights[51][6] = 3;
        layer_1_weights[52][6] = 2;
        layer_1_weights[53][6] = 1;
        layer_1_weights[54][6] = 0;
        layer_1_weights[55][6] = 1;
        layer_1_weights[56][6] = 8;
        layer_1_weights[57][6] = 11;
        layer_1_weights[58][6] = 9;
        layer_1_weights[59][6] = -20;
        layer_1_weights[60][6] = -22;
        layer_1_weights[61][6] = 3;
        layer_1_weights[62][6] = 1;
        layer_1_weights[63][6] = 1;
        layer_1_weights[64][6] = -4;
        layer_1_weights[65][6] = -4;
        layer_1_weights[66][6] = -3;
        layer_1_weights[67][6] = -2;
        layer_1_weights[68][6] = 4;
        layer_1_weights[69][6] = 5;
        layer_1_weights[70][6] = 9;
        layer_1_weights[71][6] = -31;
        layer_1_weights[72][6] = -6;
        layer_1_weights[73][6] = 1;
        layer_1_weights[74][6] = -6;
        layer_1_weights[75][6] = -3;
        layer_1_weights[76][6] = -4;
        layer_1_weights[77][6] = 5;
        layer_1_weights[78][6] = -10;
        layer_1_weights[79][6] = -7;
        layer_1_weights[80][6] = -3;
        layer_1_weights[81][6] = -4;
        layer_1_weights[82][6] = -1;
        layer_1_weights[83][6] = -7;
        layer_1_weights[84][6] = -1;
        layer_1_weights[85][6] = 0;
        layer_1_weights[86][6] = 3;
        layer_1_weights[87][6] = 2;
        layer_1_weights[88][6] = 6;
        layer_1_weights[89][6] = -1;
        layer_1_weights[90][6] = -11;
        layer_1_weights[91][6] = 0;
        layer_1_weights[92][6] = -4;
        layer_1_weights[93][6] = -9;
        layer_1_weights[94][6] = -7;
        layer_1_weights[95][6] = -16;
        layer_1_weights[96][6] = 14;
        layer_1_weights[97][6] = 2;
        layer_1_weights[98][6] = 5;
        layer_1_weights[99][6] = 6;
        layer_1_weights[100][6] = 4;
        layer_1_weights[101][6] = -3;
        layer_1_weights[102][6] = -2;
        layer_1_weights[103][6] = 2;
        layer_1_weights[104][6] = 0;
        layer_1_weights[105][6] = 5;
        layer_1_weights[106][6] = 9;
        layer_1_weights[107][6] = 8;
        layer_1_weights[108][6] = -2;
        layer_1_weights[109][6] = 5;
        layer_1_weights[110][6] = 13;
        layer_1_weights[111][6] = 6;
        layer_1_weights[112][6] = 2;
        layer_1_weights[113][6] = 5;
        layer_1_weights[114][6] = 5;
        layer_1_weights[115][6] = -1;
        layer_1_weights[116][6] = 1;
        layer_1_weights[117][6] = -1;
        layer_1_weights[118][6] = 2;
        layer_1_weights[119][6] = -6;
        layer_1_weights[120][6] = -2;
        layer_1_weights[121][6] = -6;
        layer_1_weights[122][6] = -3;
        layer_1_weights[123][6] = 2;
        layer_1_weights[124][6] = 5;
        layer_1_weights[125][6] = 5;
        layer_1_weights[126][6] = 4;
        layer_1_weights[127][6] = 4;
        layer_1_weights[128][6] = 6;
        layer_1_weights[129][6] = 10;
        layer_1_weights[130][6] = 17;
        layer_1_weights[131][6] = 11;
        layer_1_weights[132][6] = -2;
        layer_1_weights[133][6] = 6;
        layer_1_weights[134][6] = 1;
        layer_1_weights[135][6] = 6;
        layer_1_weights[136][6] = 9;
        layer_1_weights[137][6] = 12;
        layer_1_weights[138][6] = 10;
        layer_1_weights[139][6] = 16;
        layer_1_weights[140][6] = 15;
        layer_1_weights[141][6] = 5;
        layer_1_weights[142][6] = -2;
        layer_1_weights[143][6] = -3;
        layer_1_weights[0][7] = -1;
        layer_1_weights[1][7] = 1;
        layer_1_weights[2][7] = 3;
        layer_1_weights[3][7] = 7;
        layer_1_weights[4][7] = 23;
        layer_1_weights[5][7] = 0;
        layer_1_weights[6][7] = -3;
        layer_1_weights[7][7] = 14;
        layer_1_weights[8][7] = 4;
        layer_1_weights[9][7] = 8;
        layer_1_weights[10][7] = -3;
        layer_1_weights[11][7] = 3;
        layer_1_weights[12][7] = 1;
        layer_1_weights[13][7] = 1;
        layer_1_weights[14][7] = 1;
        layer_1_weights[15][7] = -5;
        layer_1_weights[16][7] = -5;
        layer_1_weights[17][7] = -5;
        layer_1_weights[18][7] = -3;
        layer_1_weights[19][7] = -2;
        layer_1_weights[20][7] = 0;
        layer_1_weights[21][7] = -2;
        layer_1_weights[22][7] = 2;
        layer_1_weights[23][7] = 7;
        layer_1_weights[24][7] = -1;
        layer_1_weights[25][7] = 3;
        layer_1_weights[26][7] = 3;
        layer_1_weights[27][7] = 1;
        layer_1_weights[28][7] = 1;
        layer_1_weights[29][7] = 2;
        layer_1_weights[30][7] = 2;
        layer_1_weights[31][7] = 0;
        layer_1_weights[32][7] = 3;
        layer_1_weights[33][7] = 2;
        layer_1_weights[34][7] = 2;
        layer_1_weights[35][7] = 3;
        layer_1_weights[36][7] = 8;
        layer_1_weights[37][7] = 7;
        layer_1_weights[38][7] = 5;
        layer_1_weights[39][7] = 6;
        layer_1_weights[40][7] = 5;
        layer_1_weights[41][7] = 3;
        layer_1_weights[42][7] = -7;
        layer_1_weights[43][7] = -3;
        layer_1_weights[44][7] = 2;
        layer_1_weights[45][7] = 4;
        layer_1_weights[46][7] = 7;
        layer_1_weights[47][7] = 3;
        layer_1_weights[48][7] = 0;
        layer_1_weights[49][7] = 9;
        layer_1_weights[50][7] = 9;
        layer_1_weights[51][7] = 9;
        layer_1_weights[52][7] = 6;
        layer_1_weights[53][7] = 2;
        layer_1_weights[54][7] = 4;
        layer_1_weights[55][7] = 5;
        layer_1_weights[56][7] = 2;
        layer_1_weights[57][7] = 5;
        layer_1_weights[58][7] = 9;
        layer_1_weights[59][7] = 18;
        layer_1_weights[60][7] = 23;
        layer_1_weights[61][7] = 9;
        layer_1_weights[62][7] = 3;
        layer_1_weights[63][7] = -4;
        layer_1_weights[64][7] = -15;
        layer_1_weights[65][7] = -10;
        layer_1_weights[66][7] = -1;
        layer_1_weights[67][7] = 1;
        layer_1_weights[68][7] = -1;
        layer_1_weights[69][7] = 4;
        layer_1_weights[70][7] = 6;
        layer_1_weights[71][7] = 19;
        layer_1_weights[72][7] = 0;
        layer_1_weights[73][7] = -25;
        layer_1_weights[74][7] = -35;
        layer_1_weights[75][7] = -22;
        layer_1_weights[76][7] = -13;
        layer_1_weights[77][7] = 7;
        layer_1_weights[78][7] = 10;
        layer_1_weights[79][7] = -5;
        layer_1_weights[80][7] = -7;
        layer_1_weights[81][7] = -6;
        layer_1_weights[82][7] = -6;
        layer_1_weights[83][7] = 7;
        layer_1_weights[84][7] = -5;
        layer_1_weights[85][7] = -36;
        layer_1_weights[86][7] = -11;
        layer_1_weights[87][7] = -2;
        layer_1_weights[88][7] = 9;
        layer_1_weights[89][7] = 15;
        layer_1_weights[90][7] = 3;
        layer_1_weights[91][7] = -6;
        layer_1_weights[92][7] = -7;
        layer_1_weights[93][7] = -3;
        layer_1_weights[94][7] = 2;
        layer_1_weights[95][7] = 11;
        layer_1_weights[96][7] = -4;
        layer_1_weights[97][7] = 2;
        layer_1_weights[98][7] = -2;
        layer_1_weights[99][7] = 6;
        layer_1_weights[100][7] = 9;
        layer_1_weights[101][7] = 7;
        layer_1_weights[102][7] = -4;
        layer_1_weights[103][7] = -3;
        layer_1_weights[104][7] = -2;
        layer_1_weights[105][7] = -4;
        layer_1_weights[106][7] = 4;
        layer_1_weights[107][7] = 5;
        layer_1_weights[108][7] = 9;
        layer_1_weights[109][7] = 0;
        layer_1_weights[110][7] = 8;
        layer_1_weights[111][7] = 1;
        layer_1_weights[112][7] = 0;
        layer_1_weights[113][7] = 5;
        layer_1_weights[114][7] = 7;
        layer_1_weights[115][7] = 6;
        layer_1_weights[116][7] = 8;
        layer_1_weights[117][7] = 4;
        layer_1_weights[118][7] = -3;
        layer_1_weights[119][7] = 2;
        layer_1_weights[120][7] = 2;
        layer_1_weights[121][7] = -12;
        layer_1_weights[122][7] = -2;
        layer_1_weights[123][7] = 1;
        layer_1_weights[124][7] = 2;
        layer_1_weights[125][7] = 6;
        layer_1_weights[126][7] = 7;
        layer_1_weights[127][7] = 4;
        layer_1_weights[128][7] = 4;
        layer_1_weights[129][7] = 0;
        layer_1_weights[130][7] = 6;
        layer_1_weights[131][7] = 15;
        layer_1_weights[132][7] = -3;
        layer_1_weights[133][7] = -9;
        layer_1_weights[134][7] = -5;
        layer_1_weights[135][7] = -3;
        layer_1_weights[136][7] = 1;
        layer_1_weights[137][7] = -2;
        layer_1_weights[138][7] = -1;
        layer_1_weights[139][7] = 1;
        layer_1_weights[140][7] = 0;
        layer_1_weights[141][7] = -1;
        layer_1_weights[142][7] = 1;
        layer_1_weights[143][7] = 2;
        layer_1_biases[0] = 2;
        layer_1_biases[1] = 5;
        layer_1_biases[2] = 5;
        layer_1_biases[3] = 4;
        layer_1_biases[4] = -22;
        layer_1_biases[5] = -1;
        layer_1_biases[6] = -13;
        layer_1_biases[7] = -14;
        layer_2_weights[0][0] = 9;
        layer_2_weights[1][0] = 3;
        layer_2_weights[2][0] = -23;
        layer_2_weights[3][0] = -12;
        layer_2_weights[4][0] = -16;
        layer_2_weights[5][0] = 11;
        layer_2_weights[6][0] = 13;
        layer_2_weights[7][0] = -12;
        layer_2_weights[0][1] = -2;
        layer_2_weights[1][1] = -28;
        layer_2_weights[2][1] = 20;
        layer_2_weights[3][1] = 7;
        layer_2_weights[4][1] = -15;
        layer_2_weights[5][1] = -8;
        layer_2_weights[6][1] = -12;
        layer_2_weights[7][1] = 10;
        layer_2_weights[0][2] = -15;
        layer_2_weights[1][2] = -8;
        layer_2_weights[2][2] = -6;
        layer_2_weights[3][2] = -17;
        layer_2_weights[4][2] = 7;
        layer_2_weights[5][2] = 15;
        layer_2_weights[6][2] = 6;
        layer_2_weights[7][2] = 26;
        layer_2_weights[0][3] = -9;
        layer_2_weights[1][3] = 8;
        layer_2_weights[2][3] = 13;
        layer_2_weights[3][3] = -9;
        layer_2_weights[4][3] = -4;
        layer_2_weights[5][3] = 5;
        layer_2_weights[6][3] = -1;
        layer_2_weights[7][3] = 6;
        layer_2_weights[0][4] = 7;
        layer_2_weights[1][4] = 5;
        layer_2_weights[2][4] = -6;
        layer_2_weights[3][4] = 0;
        layer_2_weights[4][4] = 17;
        layer_2_weights[5][4] = -11;
        layer_2_weights[6][4] = -35;
        layer_2_weights[7][4] = -12;
        layer_2_weights[0][5] = 13;
        layer_2_weights[1][5] = 1;
        layer_2_weights[2][5] = 7;
        layer_2_weights[3][5] = -28;
        layer_2_weights[4][5] = -6;
        layer_2_weights[5][5] = -6;
        layer_2_weights[6][5] = -8;
        layer_2_weights[7][5] = -4;
        layer_2_weights[0][6] = 15;
        layer_2_weights[1][6] = -20;
        layer_2_weights[2][6] = -21;
        layer_2_weights[3][6] = -2;
        layer_2_weights[4][6] = -6;
        layer_2_weights[5][6] = 18;
        layer_2_weights[6][6] = -9;
        layer_2_weights[7][6] = -6;
        layer_2_weights[0][7] = -7;
        layer_2_weights[1][7] = 16;
        layer_2_weights[2][7] = -22;
        layer_2_weights[3][7] = 10;
        layer_2_weights[4][7] = -23;
        layer_2_weights[5][7] = -5;
        layer_2_weights[6][7] = -10;
        layer_2_weights[7][7] = 9;
        layer_2_weights[0][8] = 11;
        layer_2_weights[1][8] = -1;
        layer_2_weights[2][8] = 6;
        layer_2_weights[3][8] = -9;
        layer_2_weights[4][8] = 8;
        layer_2_weights[5][8] = -3;
        layer_2_weights[6][8] = 0;
        layer_2_weights[7][8] = 11;
        layer_2_weights[0][9] = 1;
        layer_2_weights[1][9] = -1;
        layer_2_weights[2][9] = 1;
        layer_2_weights[3][9] = 10;
        layer_2_weights[4][9] = 7;
        layer_2_weights[5][9] = -26;
        layer_2_weights[6][9] = 8;
        layer_2_weights[7][9] = -27;
        layer_2_biases[0] = -11;
        layer_2_biases[1] = 14;
        layer_2_biases[2] = 20;
        layer_2_biases[3] = -23;
        layer_2_biases[4] = 4;
        layer_2_biases[5] = 47;
        layer_2_biases[6] = -12;
        layer_2_biases[7] = 19;
        layer_2_biases[8] = -55;
        layer_2_biases[9] = -6;
    end

    integer i, j, k;
    always @(*) begin
        if (predict) begin

            // Layer 1 Computation
            for (j = 0; j < 8; j = j + 1) begin
                layer_1_outputs[j] = layer_1_biases[j]; // Initialize with bias
                for (k = 0; k < 144; k = k + 1) begin
                    if (inp[k] == 1)
                        layer_1_outputs[j] = layer_1_outputs[j] + layer_1_weights[k][j];
                end
            end

            // Layer 2 Computation
            for (j = 0; j < 10; j = j + 1) begin
                layer_2_outputs[j] = layer_2_biases[j]; // Initialize with bias
                for (k = 0; k < 8; k = k + 1) begin
                    layer_2_outputs[j] = layer_2_outputs[j] + layer_1_outputs[k] * layer_2_weights[k][j];
                end
                // Apply ReLU
                if (layer_2_outputs[j] < 0)
                    layer_2_outputs[j] = 0;
            end

            // Winner-takes-all logic
            max_val = layer_2_outputs[0];
            max_idx = 0;
            for (i = 1; i < 10; i = i + 1) begin
                if (layer_2_outputs[i] > max_val) begin
                    max_val = layer_2_outputs[i];
                    max_idx = i;
                end
            end
            class = max_idx;

        end else begin
            class = 10;
        end
    end

endmodule